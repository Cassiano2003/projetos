entity mux_8_tb is
end mux_8_tb;

architecture teste of mux_8_tb is
    signal d0,d1,d2,d3,d4,d5,d6,d7,c1,c2,c3,c4,c5,r : bit;
    begin
        m : entity work.mux_8(dataflow)
            port map(d0,d1,d2,d3,d4,d5,d6,d7,c1,c2,c3,c4,c5,r);
        estimulo_checagem : process is
            type linha_tv is record
            d0,d1,d2,d3,d4,d5,d6,d7,c1,c2,c3,c4,c5, r: bit;
            end record;
            type vet_linha_tv is array (0 to 8191) of linha_tv;
            constant tabela_verdade : vet_linha_tv := 
            (
            --  d0,d1,d2,d3,d4,d5,d6,d7,c1,c2,c3,c4,c5,r
            ('0','0','0','0','0','0','0','0','0','0','0','0','0','0'),
            ('0','0','0','0','0','0','0','0','0','0','0','0','1','0'),
            ('0','0','0','0','0','0','0','0','0','0','0','1','0','0'),
            ('0','0','0','0','0','0','0','0','0','0','0','1','1','0'),
            ('0','0','0','0','0','0','0','0','0','0','1','0','0','0'),
            ('0','0','0','0','0','0','0','0','0','0','1','0','1','0'),
            ('0','0','0','0','0','0','0','0','0','0','1','1','0','0'),
            ('0','0','0','0','0','0','0','0','0','0','1','1','1','0'),
            ('0','0','0','0','0','0','0','0','0','1','0','0','0','0'),
            ('0','0','0','0','0','0','0','0','0','1','0','0','1','0'),
            ('0','0','0','0','0','0','0','0','0','1','0','1','0','0'),
            ('0','0','0','0','0','0','0','0','0','1','0','1','1','0'),
            ('0','0','0','0','0','0','0','0','0','1','1','0','0','0'),
            ('0','0','0','0','0','0','0','0','0','1','1','0','1','0'),
            ('0','0','0','0','0','0','0','0','0','1','1','1','0','0'),
            ('0','0','0','0','0','0','0','0','0','1','1','1','1','0'),
            ('0','0','0','0','0','0','0','0','1','0','0','0','0','0'),
            ('0','0','0','0','0','0','0','0','1','0','0','0','1','0'),
            ('0','0','0','0','0','0','0','0','1','0','0','1','0','0'),
            ('0','0','0','0','0','0','0','0','1','0','0','1','1','0'),
            ('0','0','0','0','0','0','0','0','1','0','1','0','0','0'),
            ('0','0','0','0','0','0','0','0','1','0','1','0','1','0'),
            ('0','0','0','0','0','0','0','0','1','0','1','1','0','0'),
            ('0','0','0','0','0','0','0','0','1','0','1','1','1','0'),
            ('0','0','0','0','0','0','0','0','1','1','0','0','0','0'),
            ('0','0','0','0','0','0','0','0','1','1','0','0','1','0'),
            ('0','0','0','0','0','0','0','0','1','1','0','1','0','0'),
            ('0','0','0','0','0','0','0','0','1','1','0','1','1','0'),
            ('0','0','0','0','0','0','0','0','1','1','1','0','0','0'),
            ('0','0','0','0','0','0','0','0','1','1','1','0','1','0'),
            ('0','0','0','0','0','0','0','0','1','1','1','1','0','0'),
            ('0','0','0','0','0','0','0','0','1','1','1','1','1','0'),
            ('0','0','0','0','0','0','0','1','0','0','0','0','0','0'),
            ('0','0','0','0','0','0','0','1','0','0','0','0','1','0'),
            ('0','0','0','0','0','0','0','1','0','0','0','1','0','0'),
            ('0','0','0','0','0','0','0','1','0','0','0','1','1','0'),
            ('0','0','0','0','0','0','0','1','0','0','1','0','0','0'),
            ('0','0','0','0','0','0','0','1','0','0','1','0','1','0'),
            ('0','0','0','0','0','0','0','1','0','0','1','1','0','0'),
            ('0','0','0','0','0','0','0','1','0','0','1','1','1','0'),
            ('0','0','0','0','0','0','0','1','0','1','0','0','0','0'),
            ('0','0','0','0','0','0','0','1','0','1','0','0','1','0'),
            ('0','0','0','0','0','0','0','1','0','1','0','1','0','0'),
            ('0','0','0','0','0','0','0','1','0','1','0','1','1','0'),
            ('0','0','0','0','0','0','0','1','0','1','1','0','0','0'),
            ('0','0','0','0','0','0','0','1','0','1','1','0','1','0'),
            ('0','0','0','0','0','0','0','1','0','1','1','1','0','0'),
            ('0','0','0','0','0','0','0','1','0','1','1','1','1','0'),
            ('0','0','0','0','0','0','0','1','1','0','0','0','0','0'),
            ('0','0','0','0','0','0','0','1','1','0','0','0','1','0'),
            ('0','0','0','0','0','0','0','1','1','0','0','1','0','0'),
            ('0','0','0','0','0','0','0','1','1','0','0','1','1','0'),
            ('0','0','0','0','0','0','0','1','1','0','1','0','0','0'),
            ('0','0','0','0','0','0','0','1','1','0','1','0','1','0'),
            ('0','0','0','0','0','0','0','1','1','0','1','1','0','0'),
            ('0','0','0','0','0','0','0','1','1','0','1','1','1','0'),
            ('0','0','0','0','0','0','0','1','1','1','0','0','0','0'),
            ('0','0','0','0','0','0','0','1','1','1','0','0','1','0'),
            ('0','0','0','0','0','0','0','1','1','1','0','1','0','0'),
            ('0','0','0','0','0','0','0','1','1','1','0','1','1','0'),
            ('0','0','0','0','0','0','0','1','1','1','1','0','0','0'),
            ('0','0','0','0','0','0','0','1','1','1','1','0','1','0'),
            ('0','0','0','0','0','0','0','1','1','1','1','1','0','0'),
            ('0','0','0','0','0','0','0','1','1','1','1','1','1','0'),
            ('0','0','0','0','0','0','1','0','0','0','0','0','0','0'),
            ('0','0','0','0','0','0','1','0','0','0','0','0','1','0'),
            ('0','0','0','0','0','0','1','0','0','0','0','1','0','0'),
            ('0','0','0','0','0','0','1','0','0','0','0','1','1','0'),
            ('0','0','0','0','0','0','1','0','0','0','1','0','0','0'),
            ('0','0','0','0','0','0','1','0','0','0','1','0','1','0'),
            ('0','0','0','0','0','0','1','0','0','0','1','1','0','0'),
            ('0','0','0','0','0','0','1','0','0','0','1','1','1','0'),
            ('0','0','0','0','0','0','1','0','0','1','0','0','0','0'),
            ('0','0','0','0','0','0','1','0','0','1','0','0','1','0'),
            ('0','0','0','0','0','0','1','0','0','1','0','1','0','0'),
            ('0','0','0','0','0','0','1','0','0','1','0','1','1','0'),
            ('0','0','0','0','0','0','1','0','0','1','1','0','0','0'),
            ('0','0','0','0','0','0','1','0','0','1','1','0','1','0'),
            ('0','0','0','0','0','0','1','0','0','1','1','1','0','0'),
            ('0','0','0','0','0','0','1','0','0','1','1','1','1','0'),
            ('0','0','0','0','0','0','1','0','1','0','0','0','0','0'),
            ('0','0','0','0','0','0','1','0','1','0','0','0','1','0'),
            ('0','0','0','0','0','0','1','0','1','0','0','1','0','0'),
            ('0','0','0','0','0','0','1','0','1','0','0','1','1','0'),
            ('0','0','0','0','0','0','1','0','1','0','1','0','0','0'),
            ('0','0','0','0','0','0','1','0','1','0','1','0','1','0'),
            ('0','0','0','0','0','0','1','0','1','0','1','1','0','0'),
            ('0','0','0','0','0','0','1','0','1','0','1','1','1','0'),
            ('0','0','0','0','0','0','1','0','1','1','0','0','0','0'),
            ('0','0','0','0','0','0','1','0','1','1','0','0','1','0'),
            ('0','0','0','0','0','0','1','0','1','1','0','1','0','0'),
            ('0','0','0','0','0','0','1','0','1','1','0','1','1','0'),
            ('0','0','0','0','0','0','1','0','1','1','1','0','0','0'),
            ('0','0','0','0','0','0','1','0','1','1','1','0','1','0'),
            ('0','0','0','0','0','0','1','0','1','1','1','1','0','0'),
            ('0','0','0','0','0','0','1','0','1','1','1','1','1','0'),
            ('0','0','0','0','0','0','1','1','0','0','0','0','0','0'),
            ('0','0','0','0','0','0','1','1','0','0','0','0','1','0'),
            ('0','0','0','0','0','0','1','1','0','0','0','1','0','0'),
            ('0','0','0','0','0','0','1','1','0','0','0','1','1','0'),
            ('0','0','0','0','0','0','1','1','0','0','1','0','0','0'),
            ('0','0','0','0','0','0','1','1','0','0','1','0','1','0'),
            ('0','0','0','0','0','0','1','1','0','0','1','1','0','0'),
            ('0','0','0','0','0','0','1','1','0','0','1','1','1','0'),
            ('0','0','0','0','0','0','1','1','0','1','0','0','0','0'),
            ('0','0','0','0','0','0','1','1','0','1','0','0','1','0'),
            ('0','0','0','0','0','0','1','1','0','1','0','1','0','0'),
            ('0','0','0','0','0','0','1','1','0','1','0','1','1','0'),
            ('0','0','0','0','0','0','1','1','0','1','1','0','0','0'),
            ('0','0','0','0','0','0','1','1','0','1','1','0','1','0'),
            ('0','0','0','0','0','0','1','1','0','1','1','1','0','0'),
            ('0','0','0','0','0','0','1','1','0','1','1','1','1','0'),
            ('0','0','0','0','0','0','1','1','1','0','0','0','0','0'),
            ('0','0','0','0','0','0','1','1','1','0','0','0','1','0'),
            ('0','0','0','0','0','0','1','1','1','0','0','1','0','0'),
            ('0','0','0','0','0','0','1','1','1','0','0','1','1','0'),
            ('0','0','0','0','0','0','1','1','1','0','1','0','0','0'),
            ('0','0','0','0','0','0','1','1','1','0','1','0','1','0'),
            ('0','0','0','0','0','0','1','1','1','0','1','1','0','0'),
            ('0','0','0','0','0','0','1','1','1','0','1','1','1','0'),
            ('0','0','0','0','0','0','1','1','1','1','0','0','0','0'),
            ('0','0','0','0','0','0','1','1','1','1','0','0','1','0'),
            ('0','0','0','0','0','0','1','1','1','1','0','1','0','0'),
            ('0','0','0','0','0','0','1','1','1','1','0','1','1','0'),
            ('0','0','0','0','0','0','1','1','1','1','1','0','0','0'),
            ('0','0','0','0','0','0','1','1','1','1','1','0','1','0'),
            ('0','0','0','0','0','0','1','1','1','1','1','1','0','0'),
            ('0','0','0','0','0','0','1','1','1','1','1','1','1','0'),
            ('0','0','0','0','0','1','0','0','0','0','0','0','0','0'),
            ('0','0','0','0','0','1','0','0','0','0','0','0','1','0'),
            ('0','0','0','0','0','1','0','0','0','0','0','1','0','0'),
            ('0','0','0','0','0','1','0','0','0','0','0','1','1','0'),
            ('0','0','0','0','0','1','0','0','0','0','1','0','0','0'),
            ('0','0','0','0','0','1','0','0','0','0','1','0','1','0'),
            ('0','0','0','0','0','1','0','0','0','0','1','1','0','0'),
            ('0','0','0','0','0','1','0','0','0','0','1','1','1','0'),
            ('0','0','0','0','0','1','0','0','0','1','0','0','0','0'),
            ('0','0','0','0','0','1','0','0','0','1','0','0','1','0'),
            ('0','0','0','0','0','1','0','0','0','1','0','1','0','0'),
            ('0','0','0','0','0','1','0','0','0','1','0','1','1','0'),
            ('0','0','0','0','0','1','0','0','0','1','1','0','0','0'),
            ('0','0','0','0','0','1','0','0','0','1','1','0','1','0'),
            ('0','0','0','0','0','1','0','0','0','1','1','1','0','0'),
            ('0','0','0','0','0','1','0','0','0','1','1','1','1','0'),
            ('0','0','0','0','0','1','0','0','1','0','0','0','0','0'),
            ('0','0','0','0','0','1','0','0','1','0','0','0','1','0'),
            ('0','0','0','0','0','1','0','0','1','0','0','1','0','0'),
            ('0','0','0','0','0','1','0','0','1','0','0','1','1','0'),
            ('0','0','0','0','0','1','0','0','1','0','1','0','0','0'),
            ('0','0','0','0','0','1','0','0','1','0','1','0','1','0'),
            ('0','0','0','0','0','1','0','0','1','0','1','1','0','0'),
            ('0','0','0','0','0','1','0','0','1','0','1','1','1','0'),
            ('0','0','0','0','0','1','0','0','1','1','0','0','0','0'),
            ('0','0','0','0','0','1','0','0','1','1','0','0','1','0'),
            ('0','0','0','0','0','1','0','0','1','1','0','1','0','0'),
            ('0','0','0','0','0','1','0','0','1','1','0','1','1','0'),
            ('0','0','0','0','0','1','0','0','1','1','1','0','0','0'),
            ('0','0','0','0','0','1','0','0','1','1','1','0','1','0'),
            ('0','0','0','0','0','1','0','0','1','1','1','1','0','0'),
            ('0','0','0','0','0','1','0','0','1','1','1','1','1','0'),
            ('0','0','0','0','0','1','0','1','0','0','0','0','0','0'),
            ('0','0','0','0','0','1','0','1','0','0','0','0','1','0'),
            ('0','0','0','0','0','1','0','1','0','0','0','1','0','0'),
            ('0','0','0','0','0','1','0','1','0','0','0','1','1','0'),
            ('0','0','0','0','0','1','0','1','0','0','1','0','0','0'),
            ('0','0','0','0','0','1','0','1','0','0','1','0','1','0'),
            ('0','0','0','0','0','1','0','1','0','0','1','1','0','0'),
            ('0','0','0','0','0','1','0','1','0','0','1','1','1','0'),
            ('0','0','0','0','0','1','0','1','0','1','0','0','0','0'),
            ('0','0','0','0','0','1','0','1','0','1','0','0','1','0'),
            ('0','0','0','0','0','1','0','1','0','1','0','1','0','0'),
            ('0','0','0','0','0','1','0','1','0','1','0','1','1','0'),
            ('0','0','0','0','0','1','0','1','0','1','1','0','0','0'),
            ('0','0','0','0','0','1','0','1','0','1','1','0','1','0'),
            ('0','0','0','0','0','1','0','1','0','1','1','1','0','0'),
            ('0','0','0','0','0','1','0','1','0','1','1','1','1','0'),
            ('0','0','0','0','0','1','0','1','1','0','0','0','0','0'),
            ('0','0','0','0','0','1','0','1','1','0','0','0','1','0'),
            ('0','0','0','0','0','1','0','1','1','0','0','1','0','0'),
            ('0','0','0','0','0','1','0','1','1','0','0','1','1','0'),
            ('0','0','0','0','0','1','0','1','1','0','1','0','0','0'),
            ('0','0','0','0','0','1','0','1','1','0','1','0','1','0'),
            ('0','0','0','0','0','1','0','1','1','0','1','1','0','0'),
            ('0','0','0','0','0','1','0','1','1','0','1','1','1','0'),
            ('0','0','0','0','0','1','0','1','1','1','0','0','0','0'),
            ('0','0','0','0','0','1','0','1','1','1','0','0','1','0'),
            ('0','0','0','0','0','1','0','1','1','1','0','1','0','0'),
            ('0','0','0','0','0','1','0','1','1','1','0','1','1','0'),
            ('0','0','0','0','0','1','0','1','1','1','1','0','0','0'),
            ('0','0','0','0','0','1','0','1','1','1','1','0','1','0'),
            ('0','0','0','0','0','1','0','1','1','1','1','1','0','0'),
            ('0','0','0','0','0','1','0','1','1','1','1','1','1','0'),
            ('0','0','0','0','0','1','1','0','0','0','0','0','0','0'),
            ('0','0','0','0','0','1','1','0','0','0','0','0','1','0'),
            ('0','0','0','0','0','1','1','0','0','0','0','1','0','0'),
            ('0','0','0','0','0','1','1','0','0','0','0','1','1','0'),
            ('0','0','0','0','0','1','1','0','0','0','1','0','0','0'),
            ('0','0','0','0','0','1','1','0','0','0','1','0','1','0'),
            ('0','0','0','0','0','1','1','0','0','0','1','1','0','0'),
            ('0','0','0','0','0','1','1','0','0','0','1','1','1','0'),
            ('0','0','0','0','0','1','1','0','0','1','0','0','0','0'),
            ('0','0','0','0','0','1','1','0','0','1','0','0','1','0'),
            ('0','0','0','0','0','1','1','0','0','1','0','1','0','0'),
            ('0','0','0','0','0','1','1','0','0','1','0','1','1','0'),
            ('0','0','0','0','0','1','1','0','0','1','1','0','0','0'),
            ('0','0','0','0','0','1','1','0','0','1','1','0','1','0'),
            ('0','0','0','0','0','1','1','0','0','1','1','1','0','0'),
            ('0','0','0','0','0','1','1','0','0','1','1','1','1','0'),
            ('0','0','0','0','0','1','1','0','1','0','0','0','0','0'),
            ('0','0','0','0','0','1','1','0','1','0','0','0','1','0'),
            ('0','0','0','0','0','1','1','0','1','0','0','1','0','0'),
            ('0','0','0','0','0','1','1','0','1','0','0','1','1','0'),
            ('0','0','0','0','0','1','1','0','1','0','1','0','0','0'),
            ('0','0','0','0','0','1','1','0','1','0','1','0','1','0'),
            ('0','0','0','0','0','1','1','0','1','0','1','1','0','0'),
            ('0','0','0','0','0','1','1','0','1','0','1','1','1','0'),
            ('0','0','0','0','0','1','1','0','1','1','0','0','0','0'),
            ('0','0','0','0','0','1','1','0','1','1','0','0','1','0'),
            ('0','0','0','0','0','1','1','0','1','1','0','1','0','0'),
            ('0','0','0','0','0','1','1','0','1','1','0','1','1','0'),
            ('0','0','0','0','0','1','1','0','1','1','1','0','0','0'),
            ('0','0','0','0','0','1','1','0','1','1','1','0','1','0'),
            ('0','0','0','0','0','1','1','0','1','1','1','1','0','0'),
            ('0','0','0','0','0','1','1','0','1','1','1','1','1','0'),
            ('0','0','0','0','0','1','1','1','0','0','0','0','0','0'),
            ('0','0','0','0','0','1','1','1','0','0','0','0','1','0'),
            ('0','0','0','0','0','1','1','1','0','0','0','1','0','0'),
            ('0','0','0','0','0','1','1','1','0','0','0','1','1','0'),
            ('0','0','0','0','0','1','1','1','0','0','1','0','0','0'),
            ('0','0','0','0','0','1','1','1','0','0','1','0','1','0'),
            ('0','0','0','0','0','1','1','1','0','0','1','1','0','0'),
            ('0','0','0','0','0','1','1','1','0','0','1','1','1','0'),
            ('0','0','0','0','0','1','1','1','0','1','0','0','0','0'),
            ('0','0','0','0','0','1','1','1','0','1','0','0','1','0'),
            ('0','0','0','0','0','1','1','1','0','1','0','1','0','0'),
            ('0','0','0','0','0','1','1','1','0','1','0','1','1','0'),
            ('0','0','0','0','0','1','1','1','0','1','1','0','0','0'),
            ('0','0','0','0','0','1','1','1','0','1','1','0','1','0'),
            ('0','0','0','0','0','1','1','1','0','1','1','1','0','0'),
            ('0','0','0','0','0','1','1','1','0','1','1','1','1','0'),
            ('0','0','0','0','0','1','1','1','1','0','0','0','0','0'),
            ('0','0','0','0','0','1','1','1','1','0','0','0','1','0'),
            ('0','0','0','0','0','1','1','1','1','0','0','1','0','0'),
            ('0','0','0','0','0','1','1','1','1','0','0','1','1','0'),
            ('0','0','0','0','0','1','1','1','1','0','1','0','0','0'),
            ('0','0','0','0','0','1','1','1','1','0','1','0','1','0'),
            ('0','0','0','0','0','1','1','1','1','0','1','1','0','0'),
            ('0','0','0','0','0','1','1','1','1','0','1','1','1','0'),
            ('0','0','0','0','0','1','1','1','1','1','0','0','0','0'),
            ('0','0','0','0','0','1','1','1','1','1','0','0','1','0'),
            ('0','0','0','0','0','1','1','1','1','1','0','1','0','0'),
            ('0','0','0','0','0','1','1','1','1','1','0','1','1','0'),
            ('0','0','0','0','0','1','1','1','1','1','1','0','0','0'),
            ('0','0','0','0','0','1','1','1','1','1','1','0','1','0'),
            ('0','0','0','0','0','1','1','1','1','1','1','1','0','0'),
            ('0','0','0','0','0','1','1','1','1','1','1','1','1','0'),
            ('0','0','0','0','1','0','0','0','0','0','0','0','0','0'),
            ('0','0','0','0','1','0','0','0','0','0','0','0','1','0'),
            ('0','0','0','0','1','0','0','0','0','0','0','1','0','0'),
            ('0','0','0','0','1','0','0','0','0','0','0','1','1','0'),
            ('0','0','0','0','1','0','0','0','0','0','1','0','0','0'),
            ('0','0','0','0','1','0','0','0','0','0','1','0','1','0'),
            ('0','0','0','0','1','0','0','0','0','0','1','1','0','0'),
            ('0','0','0','0','1','0','0','0','0','0','1','1','1','0'),
            ('0','0','0','0','1','0','0','0','0','1','0','0','0','0'),
            ('0','0','0','0','1','0','0','0','0','1','0','0','1','0'),
            ('0','0','0','0','1','0','0','0','0','1','0','1','0','0'),
            ('0','0','0','0','1','0','0','0','0','1','0','1','1','0'),
            ('0','0','0','0','1','0','0','0','0','1','1','0','0','0'),
            ('0','0','0','0','1','0','0','0','0','1','1','0','1','0'),
            ('0','0','0','0','1','0','0','0','0','1','1','1','0','0'),
            ('0','0','0','0','1','0','0','0','0','1','1','1','1','0'),
            ('0','0','0','0','1','0','0','0','1','0','0','0','0','0'),
            ('0','0','0','0','1','0','0','0','1','0','0','0','1','0'),
            ('0','0','0','0','1','0','0','0','1','0','0','1','0','0'),
            ('0','0','0','0','1','0','0','0','1','0','0','1','1','0'),
            ('0','0','0','0','1','0','0','0','1','0','1','0','0','0'),
            ('0','0','0','0','1','0','0','0','1','0','1','0','1','0'),
            ('0','0','0','0','1','0','0','0','1','0','1','1','0','0'),
            ('0','0','0','0','1','0','0','0','1','0','1','1','1','0'),
            ('0','0','0','0','1','0','0','0','1','1','0','0','0','0'),
            ('0','0','0','0','1','0','0','0','1','1','0','0','1','0'),
            ('0','0','0','0','1','0','0','0','1','1','0','1','0','0'),
            ('0','0','0','0','1','0','0','0','1','1','0','1','1','0'),
            ('0','0','0','0','1','0','0','0','1','1','1','0','0','0'),
            ('0','0','0','0','1','0','0','0','1','1','1','0','1','0'),
            ('0','0','0','0','1','0','0','0','1','1','1','1','0','0'),
            ('0','0','0','0','1','0','0','0','1','1','1','1','1','0'),
            ('0','0','0','0','1','0','0','1','0','0','0','0','0','0'),
            ('0','0','0','0','1','0','0','1','0','0','0','0','1','0'),
            ('0','0','0','0','1','0','0','1','0','0','0','1','0','0'),
            ('0','0','0','0','1','0','0','1','0','0','0','1','1','0'),
            ('0','0','0','0','1','0','0','1','0','0','1','0','0','0'),
            ('0','0','0','0','1','0','0','1','0','0','1','0','1','0'),
            ('0','0','0','0','1','0','0','1','0','0','1','1','0','0'),
            ('0','0','0','0','1','0','0','1','0','0','1','1','1','0'),
            ('0','0','0','0','1','0','0','1','0','1','0','0','0','0'),
            ('0','0','0','0','1','0','0','1','0','1','0','0','1','0'),
            ('0','0','0','0','1','0','0','1','0','1','0','1','0','0'),
            ('0','0','0','0','1','0','0','1','0','1','0','1','1','0'),
            ('0','0','0','0','1','0','0','1','0','1','1','0','0','0'),
            ('0','0','0','0','1','0','0','1','0','1','1','0','1','0'),
            ('0','0','0','0','1','0','0','1','0','1','1','1','0','0'),
            ('0','0','0','0','1','0','0','1','0','1','1','1','1','0'),
            ('0','0','0','0','1','0','0','1','1','0','0','0','0','0'),
            ('0','0','0','0','1','0','0','1','1','0','0','0','1','0'),
            ('0','0','0','0','1','0','0','1','1','0','0','1','0','0'),
            ('0','0','0','0','1','0','0','1','1','0','0','1','1','0'),
            ('0','0','0','0','1','0','0','1','1','0','1','0','0','0'),
            ('0','0','0','0','1','0','0','1','1','0','1','0','1','0'),
            ('0','0','0','0','1','0','0','1','1','0','1','1','0','0'),
            ('0','0','0','0','1','0','0','1','1','0','1','1','1','0'),
            ('0','0','0','0','1','0','0','1','1','1','0','0','0','0'),
            ('0','0','0','0','1','0','0','1','1','1','0','0','1','0'),
            ('0','0','0','0','1','0','0','1','1','1','0','1','0','0'),
            ('0','0','0','0','1','0','0','1','1','1','0','1','1','0'),
            ('0','0','0','0','1','0','0','1','1','1','1','0','0','0'),
            ('0','0','0','0','1','0','0','1','1','1','1','0','1','0'),
            ('0','0','0','0','1','0','0','1','1','1','1','1','0','0'),
            ('0','0','0','0','1','0','0','1','1','1','1','1','1','0'),
            ('0','0','0','0','1','0','1','0','0','0','0','0','0','0'),
            ('0','0','0','0','1','0','1','0','0','0','0','0','1','0'),
            ('0','0','0','0','1','0','1','0','0','0','0','1','0','0'),
            ('0','0','0','0','1','0','1','0','0','0','0','1','1','0'),
            ('0','0','0','0','1','0','1','0','0','0','1','0','0','0'),
            ('0','0','0','0','1','0','1','0','0','0','1','0','1','0'),
            ('0','0','0','0','1','0','1','0','0','0','1','1','0','0'),
            ('0','0','0','0','1','0','1','0','0','0','1','1','1','0'),
            ('0','0','0','0','1','0','1','0','0','1','0','0','0','0'),
            ('0','0','0','0','1','0','1','0','0','1','0','0','1','0'),
            ('0','0','0','0','1','0','1','0','0','1','0','1','0','0'),
            ('0','0','0','0','1','0','1','0','0','1','0','1','1','0'),
            ('0','0','0','0','1','0','1','0','0','1','1','0','0','0'),
            ('0','0','0','0','1','0','1','0','0','1','1','0','1','0'),
            ('0','0','0','0','1','0','1','0','0','1','1','1','0','0'),
            ('0','0','0','0','1','0','1','0','0','1','1','1','1','0'),
            ('0','0','0','0','1','0','1','0','1','0','0','0','0','0'),
            ('0','0','0','0','1','0','1','0','1','0','0','0','1','0'),
            ('0','0','0','0','1','0','1','0','1','0','0','1','0','0'),
            ('0','0','0','0','1','0','1','0','1','0','0','1','1','0'),
            ('0','0','0','0','1','0','1','0','1','0','1','0','0','0'),
            ('0','0','0','0','1','0','1','0','1','0','1','0','1','0'),
            ('0','0','0','0','1','0','1','0','1','0','1','1','0','0'),
            ('0','0','0','0','1','0','1','0','1','0','1','1','1','0'),
            ('0','0','0','0','1','0','1','0','1','1','0','0','0','0'),
            ('0','0','0','0','1','0','1','0','1','1','0','0','1','0'),
            ('0','0','0','0','1','0','1','0','1','1','0','1','0','0'),
            ('0','0','0','0','1','0','1','0','1','1','0','1','1','0'),
            ('0','0','0','0','1','0','1','0','1','1','1','0','0','0'),
            ('0','0','0','0','1','0','1','0','1','1','1','0','1','0'),
            ('0','0','0','0','1','0','1','0','1','1','1','1','0','0'),
            ('0','0','0','0','1','0','1','0','1','1','1','1','1','0'),
            ('0','0','0','0','1','0','1','1','0','0','0','0','0','0'),
            ('0','0','0','0','1','0','1','1','0','0','0','0','1','0'),
            ('0','0','0','0','1','0','1','1','0','0','0','1','0','0'),
            ('0','0','0','0','1','0','1','1','0','0','0','1','1','0'),
            ('0','0','0','0','1','0','1','1','0','0','1','0','0','0'),
            ('0','0','0','0','1','0','1','1','0','0','1','0','1','0'),
            ('0','0','0','0','1','0','1','1','0','0','1','1','0','0'),
            ('0','0','0','0','1','0','1','1','0','0','1','1','1','0'),
            ('0','0','0','0','1','0','1','1','0','1','0','0','0','0'),
            ('0','0','0','0','1','0','1','1','0','1','0','0','1','0'),
            ('0','0','0','0','1','0','1','1','0','1','0','1','0','0'),
            ('0','0','0','0','1','0','1','1','0','1','0','1','1','0'),
            ('0','0','0','0','1','0','1','1','0','1','1','0','0','0'),
            ('0','0','0','0','1','0','1','1','0','1','1','0','1','0'),
            ('0','0','0','0','1','0','1','1','0','1','1','1','0','0'),
            ('0','0','0','0','1','0','1','1','0','1','1','1','1','0'),
            ('0','0','0','0','1','0','1','1','1','0','0','0','0','0'),
            ('0','0','0','0','1','0','1','1','1','0','0','0','1','0'),
            ('0','0','0','0','1','0','1','1','1','0','0','1','0','0'),
            ('0','0','0','0','1','0','1','1','1','0','0','1','1','0'),
            ('0','0','0','0','1','0','1','1','1','0','1','0','0','0'),
            ('0','0','0','0','1','0','1','1','1','0','1','0','1','0'),
            ('0','0','0','0','1','0','1','1','1','0','1','1','0','0'),
            ('0','0','0','0','1','0','1','1','1','0','1','1','1','0'),
            ('0','0','0','0','1','0','1','1','1','1','0','0','0','0'),
            ('0','0','0','0','1','0','1','1','1','1','0','0','1','0'),
            ('0','0','0','0','1','0','1','1','1','1','0','1','0','0'),
            ('0','0','0','0','1','0','1','1','1','1','0','1','1','0'),
            ('0','0','0','0','1','0','1','1','1','1','1','0','0','0'),
            ('0','0','0','0','1','0','1','1','1','1','1','0','1','0'),
            ('0','0','0','0','1','0','1','1','1','1','1','1','0','0'),
            ('0','0','0','0','1','0','1','1','1','1','1','1','1','0'),
            ('0','0','0','0','1','1','0','0','0','0','0','0','0','0'),
            ('0','0','0','0','1','1','0','0','0','0','0','0','1','0'),
            ('0','0','0','0','1','1','0','0','0','0','0','1','0','0'),
            ('0','0','0','0','1','1','0','0','0','0','0','1','1','0'),
            ('0','0','0','0','1','1','0','0','0','0','1','0','0','0'),
            ('0','0','0','0','1','1','0','0','0','0','1','0','1','0'),
            ('0','0','0','0','1','1','0','0','0','0','1','1','0','0'),
            ('0','0','0','0','1','1','0','0','0','0','1','1','1','0'),
            ('0','0','0','0','1','1','0','0','0','1','0','0','0','0'),
            ('0','0','0','0','1','1','0','0','0','1','0','0','1','0'),
            ('0','0','0','0','1','1','0','0','0','1','0','1','0','0'),
            ('0','0','0','0','1','1','0','0','0','1','0','1','1','0'),
            ('0','0','0','0','1','1','0','0','0','1','1','0','0','0'),
            ('0','0','0','0','1','1','0','0','0','1','1','0','1','0'),
            ('0','0','0','0','1','1','0','0','0','1','1','1','0','0'),
            ('0','0','0','0','1','1','0','0','0','1','1','1','1','0'),
            ('0','0','0','0','1','1','0','0','1','0','0','0','0','0'),
            ('0','0','0','0','1','1','0','0','1','0','0','0','1','0'),
            ('0','0','0','0','1','1','0','0','1','0','0','1','0','0'),
            ('0','0','0','0','1','1','0','0','1','0','0','1','1','0'),
            ('0','0','0','0','1','1','0','0','1','0','1','0','0','0'),
            ('0','0','0','0','1','1','0','0','1','0','1','0','1','0'),
            ('0','0','0','0','1','1','0','0','1','0','1','1','0','0'),
            ('0','0','0','0','1','1','0','0','1','0','1','1','1','0'),
            ('0','0','0','0','1','1','0','0','1','1','0','0','0','0'),
            ('0','0','0','0','1','1','0','0','1','1','0','0','1','0'),
            ('0','0','0','0','1','1','0','0','1','1','0','1','0','0'),
            ('0','0','0','0','1','1','0','0','1','1','0','1','1','0'),
            ('0','0','0','0','1','1','0','0','1','1','1','0','0','0'),
            ('0','0','0','0','1','1','0','0','1','1','1','0','1','0'),
            ('0','0','0','0','1','1','0','0','1','1','1','1','0','0'),
            ('0','0','0','0','1','1','0','0','1','1','1','1','1','0'),
            ('0','0','0','0','1','1','0','1','0','0','0','0','0','0'),
            ('0','0','0','0','1','1','0','1','0','0','0','0','1','0'),
            ('0','0','0','0','1','1','0','1','0','0','0','1','0','0'),
            ('0','0','0','0','1','1','0','1','0','0','0','1','1','0'),
            ('0','0','0','0','1','1','0','1','0','0','1','0','0','0'),
            ('0','0','0','0','1','1','0','1','0','0','1','0','1','0'),
            ('0','0','0','0','1','1','0','1','0','0','1','1','0','0'),
            ('0','0','0','0','1','1','0','1','0','0','1','1','1','0'),
            ('0','0','0','0','1','1','0','1','0','1','0','0','0','0'),
            ('0','0','0','0','1','1','0','1','0','1','0','0','1','0'),
            ('0','0','0','0','1','1','0','1','0','1','0','1','0','0'),
            ('0','0','0','0','1','1','0','1','0','1','0','1','1','0'),
            ('0','0','0','0','1','1','0','1','0','1','1','0','0','0'),
            ('0','0','0','0','1','1','0','1','0','1','1','0','1','0'),
            ('0','0','0','0','1','1','0','1','0','1','1','1','0','0'),
            ('0','0','0','0','1','1','0','1','0','1','1','1','1','0'),
            ('0','0','0','0','1','1','0','1','1','0','0','0','0','0'),
            ('0','0','0','0','1','1','0','1','1','0','0','0','1','0'),
            ('0','0','0','0','1','1','0','1','1','0','0','1','0','0'),
            ('0','0','0','0','1','1','0','1','1','0','0','1','1','0'),
            ('0','0','0','0','1','1','0','1','1','0','1','0','0','0'),
            ('0','0','0','0','1','1','0','1','1','0','1','0','1','0'),
            ('0','0','0','0','1','1','0','1','1','0','1','1','0','0'),
            ('0','0','0','0','1','1','0','1','1','0','1','1','1','0'),
            ('0','0','0','0','1','1','0','1','1','1','0','0','0','0'),
            ('0','0','0','0','1','1','0','1','1','1','0','0','1','0'),
            ('0','0','0','0','1','1','0','1','1','1','0','1','0','0'),
            ('0','0','0','0','1','1','0','1','1','1','0','1','1','0'),
            ('0','0','0','0','1','1','0','1','1','1','1','0','0','0'),
            ('0','0','0','0','1','1','0','1','1','1','1','0','1','0'),
            ('0','0','0','0','1','1','0','1','1','1','1','1','0','0'),
            ('0','0','0','0','1','1','0','1','1','1','1','1','1','0'),
            ('0','0','0','0','1','1','1','0','0','0','0','0','0','0'),
            ('0','0','0','0','1','1','1','0','0','0','0','0','1','0'),
            ('0','0','0','0','1','1','1','0','0','0','0','1','0','0'),
            ('0','0','0','0','1','1','1','0','0','0','0','1','1','0'),
            ('0','0','0','0','1','1','1','0','0','0','1','0','0','0'),
            ('0','0','0','0','1','1','1','0','0','0','1','0','1','0'),
            ('0','0','0','0','1','1','1','0','0','0','1','1','0','0'),
            ('0','0','0','0','1','1','1','0','0','0','1','1','1','0'),
            ('0','0','0','0','1','1','1','0','0','1','0','0','0','0'),
            ('0','0','0','0','1','1','1','0','0','1','0','0','1','0'),
            ('0','0','0','0','1','1','1','0','0','1','0','1','0','0'),
            ('0','0','0','0','1','1','1','0','0','1','0','1','1','0'),
            ('0','0','0','0','1','1','1','0','0','1','1','0','0','0'),
            ('0','0','0','0','1','1','1','0','0','1','1','0','1','0'),
            ('0','0','0','0','1','1','1','0','0','1','1','1','0','0'),
            ('0','0','0','0','1','1','1','0','0','1','1','1','1','0'),
            ('0','0','0','0','1','1','1','0','1','0','0','0','0','0'),
            ('0','0','0','0','1','1','1','0','1','0','0','0','1','0'),
            ('0','0','0','0','1','1','1','0','1','0','0','1','0','0'),
            ('0','0','0','0','1','1','1','0','1','0','0','1','1','0'),
            ('0','0','0','0','1','1','1','0','1','0','1','0','0','0'),
            ('0','0','0','0','1','1','1','0','1','0','1','0','1','0'),
            ('0','0','0','0','1','1','1','0','1','0','1','1','0','0'),
            ('0','0','0','0','1','1','1','0','1','0','1','1','1','0'),
            ('0','0','0','0','1','1','1','0','1','1','0','0','0','0'),
            ('0','0','0','0','1','1','1','0','1','1','0','0','1','0'),
            ('0','0','0','0','1','1','1','0','1','1','0','1','0','0'),
            ('0','0','0','0','1','1','1','0','1','1','0','1','1','0'),
            ('0','0','0','0','1','1','1','0','1','1','1','0','0','0'),
            ('0','0','0','0','1','1','1','0','1','1','1','0','1','0'),
            ('0','0','0','0','1','1','1','0','1','1','1','1','0','0'),
            ('0','0','0','0','1','1','1','0','1','1','1','1','1','0'),
            ('0','0','0','0','1','1','1','1','0','0','0','0','0','0'),
            ('0','0','0','0','1','1','1','1','0','0','0','0','1','0'),
            ('0','0','0','0','1','1','1','1','0','0','0','1','0','0'),
            ('0','0','0','0','1','1','1','1','0','0','0','1','1','0'),
            ('0','0','0','0','1','1','1','1','0','0','1','0','0','0'),
            ('0','0','0','0','1','1','1','1','0','0','1','0','1','0'),
            ('0','0','0','0','1','1','1','1','0','0','1','1','0','0'),
            ('0','0','0','0','1','1','1','1','0','0','1','1','1','0'),
            ('0','0','0','0','1','1','1','1','0','1','0','0','0','0'),
            ('0','0','0','0','1','1','1','1','0','1','0','0','1','0'),
            ('0','0','0','0','1','1','1','1','0','1','0','1','0','0'),
            ('0','0','0','0','1','1','1','1','0','1','0','1','1','0'),
            ('0','0','0','0','1','1','1','1','0','1','1','0','0','0'),
            ('0','0','0','0','1','1','1','1','0','1','1','0','1','0'),
            ('0','0','0','0','1','1','1','1','0','1','1','1','0','0'),
            ('0','0','0','0','1','1','1','1','0','1','1','1','1','0'),
            ('0','0','0','0','1','1','1','1','1','0','0','0','0','0'),
            ('0','0','0','0','1','1','1','1','1','0','0','0','1','0'),
            ('0','0','0','0','1','1','1','1','1','0','0','1','0','0'),
            ('0','0','0','0','1','1','1','1','1','0','0','1','1','0'),
            ('0','0','0','0','1','1','1','1','1','0','1','0','0','0'),
            ('0','0','0','0','1','1','1','1','1','0','1','0','1','0'),
            ('0','0','0','0','1','1','1','1','1','0','1','1','0','0'),
            ('0','0','0','0','1','1','1','1','1','0','1','1','1','0'),
            ('0','0','0','0','1','1','1','1','1','1','0','0','0','0'),
            ('0','0','0','0','1','1','1','1','1','1','0','0','1','0'),
            ('0','0','0','0','1','1','1','1','1','1','0','1','0','0'),
            ('0','0','0','0','1','1','1','1','1','1','0','1','1','0'),
            ('0','0','0','0','1','1','1','1','1','1','1','0','0','0'),
            ('0','0','0','0','1','1','1','1','1','1','1','0','1','0'),
            ('0','0','0','0','1','1','1','1','1','1','1','1','0','0'),
            ('0','0','0','0','1','1','1','1','1','1','1','1','1','0'),
            ('0','0','0','1','0','0','0','0','0','0','0','0','0','0'),
            ('0','0','0','1','0','0','0','0','0','0','0','0','1','0'),
            ('0','0','0','1','0','0','0','0','0','0','0','1','0','0'),
            ('0','0','0','1','0','0','0','0','0','0','0','1','1','0'),
            ('0','0','0','1','0','0','0','0','0','0','1','0','0','0'),
            ('0','0','0','1','0','0','0','0','0','0','1','0','1','0'),
            ('0','0','0','1','0','0','0','0','0','0','1','1','0','0'),
            ('0','0','0','1','0','0','0','0','0','0','1','1','1','0'),
            ('0','0','0','1','0','0','0','0','0','1','0','0','0','0'),
            ('0','0','0','1','0','0','0','0','0','1','0','0','1','0'),
            ('0','0','0','1','0','0','0','0','0','1','0','1','0','0'),
            ('0','0','0','1','0','0','0','0','0','1','0','1','1','0'),
            ('0','0','0','1','0','0','0','0','0','1','1','0','0','0'),
            ('0','0','0','1','0','0','0','0','0','1','1','0','1','0'),
            ('0','0','0','1','0','0','0','0','0','1','1','1','0','0'),
            ('0','0','0','1','0','0','0','0','0','1','1','1','1','0'),
            ('0','0','0','1','0','0','0','0','1','0','0','0','0','0'),
            ('0','0','0','1','0','0','0','0','1','0','0','0','1','0'),
            ('0','0','0','1','0','0','0','0','1','0','0','1','0','0'),
            ('0','0','0','1','0','0','0','0','1','0','0','1','1','0'),
            ('0','0','0','1','0','0','0','0','1','0','1','0','0','0'),
            ('0','0','0','1','0','0','0','0','1','0','1','0','1','0'),
            ('0','0','0','1','0','0','0','0','1','0','1','1','0','0'),
            ('0','0','0','1','0','0','0','0','1','0','1','1','1','0'),
            ('0','0','0','1','0','0','0','0','1','1','0','0','0','0'),
            ('0','0','0','1','0','0','0','0','1','1','0','0','1','0'),
            ('0','0','0','1','0','0','0','0','1','1','0','1','0','0'),
            ('0','0','0','1','0','0','0','0','1','1','0','1','1','0'),
            ('0','0','0','1','0','0','0','0','1','1','1','0','0','0'),
            ('0','0','0','1','0','0','0','0','1','1','1','0','1','0'),
            ('0','0','0','1','0','0','0','0','1','1','1','1','0','0'),
            ('0','0','0','1','0','0','0','0','1','1','1','1','1','0'),
            ('0','0','0','1','0','0','0','1','0','0','0','0','0','0'),
            ('0','0','0','1','0','0','0','1','0','0','0','0','1','0'),
            ('0','0','0','1','0','0','0','1','0','0','0','1','0','0'),
            ('0','0','0','1','0','0','0','1','0','0','0','1','1','0'),
            ('0','0','0','1','0','0','0','1','0','0','1','0','0','0'),
            ('0','0','0','1','0','0','0','1','0','0','1','0','1','0'),
            ('0','0','0','1','0','0','0','1','0','0','1','1','0','0'),
            ('0','0','0','1','0','0','0','1','0','0','1','1','1','0'),
            ('0','0','0','1','0','0','0','1','0','1','0','0','0','0'),
            ('0','0','0','1','0','0','0','1','0','1','0','0','1','0'),
            ('0','0','0','1','0','0','0','1','0','1','0','1','0','0'),
            ('0','0','0','1','0','0','0','1','0','1','0','1','1','0'),
            ('0','0','0','1','0','0','0','1','0','1','1','0','0','0'),
            ('0','0','0','1','0','0','0','1','0','1','1','0','1','0'),
            ('0','0','0','1','0','0','0','1','0','1','1','1','0','0'),
            ('0','0','0','1','0','0','0','1','0','1','1','1','1','0'),
            ('0','0','0','1','0','0','0','1','1','0','0','0','0','0'),
            ('0','0','0','1','0','0','0','1','1','0','0','0','1','0'),
            ('0','0','0','1','0','0','0','1','1','0','0','1','0','0'),
            ('0','0','0','1','0','0','0','1','1','0','0','1','1','0'),
            ('0','0','0','1','0','0','0','1','1','0','1','0','0','0'),
            ('0','0','0','1','0','0','0','1','1','0','1','0','1','0'),
            ('0','0','0','1','0','0','0','1','1','0','1','1','0','0'),
            ('0','0','0','1','0','0','0','1','1','0','1','1','1','0'),
            ('0','0','0','1','0','0','0','1','1','1','0','0','0','0'),
            ('0','0','0','1','0','0','0','1','1','1','0','0','1','0'),
            ('0','0','0','1','0','0','0','1','1','1','0','1','0','0'),
            ('0','0','0','1','0','0','0','1','1','1','0','1','1','0'),
            ('0','0','0','1','0','0','0','1','1','1','1','0','0','0'),
            ('0','0','0','1','0','0','0','1','1','1','1','0','1','0'),
            ('0','0','0','1','0','0','0','1','1','1','1','1','0','0'),
            ('0','0','0','1','0','0','0','1','1','1','1','1','1','0'),
            ('0','0','0','1','0','0','1','0','0','0','0','0','0','0'),
            ('0','0','0','1','0','0','1','0','0','0','0','0','1','0'),
            ('0','0','0','1','0','0','1','0','0','0','0','1','0','0'),
            ('0','0','0','1','0','0','1','0','0','0','0','1','1','0'),
            ('0','0','0','1','0','0','1','0','0','0','1','0','0','0'),
            ('0','0','0','1','0','0','1','0','0','0','1','0','1','0'),
            ('0','0','0','1','0','0','1','0','0','0','1','1','0','0'),
            ('0','0','0','1','0','0','1','0','0','0','1','1','1','0'),
            ('0','0','0','1','0','0','1','0','0','1','0','0','0','0'),
            ('0','0','0','1','0','0','1','0','0','1','0','0','1','0'),
            ('0','0','0','1','0','0','1','0','0','1','0','1','0','0'),
            ('0','0','0','1','0','0','1','0','0','1','0','1','1','0'),
            ('0','0','0','1','0','0','1','0','0','1','1','0','0','0'),
            ('0','0','0','1','0','0','1','0','0','1','1','0','1','0'),
            ('0','0','0','1','0','0','1','0','0','1','1','1','0','0'),
            ('0','0','0','1','0','0','1','0','0','1','1','1','1','0'),
            ('0','0','0','1','0','0','1','0','1','0','0','0','0','0'),
            ('0','0','0','1','0','0','1','0','1','0','0','0','1','0'),
            ('0','0','0','1','0','0','1','0','1','0','0','1','0','0'),
            ('0','0','0','1','0','0','1','0','1','0','0','1','1','0'),
            ('0','0','0','1','0','0','1','0','1','0','1','0','0','0'),
            ('0','0','0','1','0','0','1','0','1','0','1','0','1','0'),
            ('0','0','0','1','0','0','1','0','1','0','1','1','0','0'),
            ('0','0','0','1','0','0','1','0','1','0','1','1','1','0'),
            ('0','0','0','1','0','0','1','0','1','1','0','0','0','0'),
            ('0','0','0','1','0','0','1','0','1','1','0','0','1','0'),
            ('0','0','0','1','0','0','1','0','1','1','0','1','0','0'),
            ('0','0','0','1','0','0','1','0','1','1','0','1','1','0'),
            ('0','0','0','1','0','0','1','0','1','1','1','0','0','0'),
            ('0','0','0','1','0','0','1','0','1','1','1','0','1','0'),
            ('0','0','0','1','0','0','1','0','1','1','1','1','0','0'),
            ('0','0','0','1','0','0','1','0','1','1','1','1','1','0'),
            ('0','0','0','1','0','0','1','1','0','0','0','0','0','0'),
            ('0','0','0','1','0','0','1','1','0','0','0','0','1','0'),
            ('0','0','0','1','0','0','1','1','0','0','0','1','0','0'),
            ('0','0','0','1','0','0','1','1','0','0','0','1','1','0'),
            ('0','0','0','1','0','0','1','1','0','0','1','0','0','0'),
            ('0','0','0','1','0','0','1','1','0','0','1','0','1','0'),
            ('0','0','0','1','0','0','1','1','0','0','1','1','0','0'),
            ('0','0','0','1','0','0','1','1','0','0','1','1','1','0'),
            ('0','0','0','1','0','0','1','1','0','1','0','0','0','0'),
            ('0','0','0','1','0','0','1','1','0','1','0','0','1','0'),
            ('0','0','0','1','0','0','1','1','0','1','0','1','0','0'),
            ('0','0','0','1','0','0','1','1','0','1','0','1','1','0'),
            ('0','0','0','1','0','0','1','1','0','1','1','0','0','0'),
            ('0','0','0','1','0','0','1','1','0','1','1','0','1','0'),
            ('0','0','0','1','0','0','1','1','0','1','1','1','0','0'),
            ('0','0','0','1','0','0','1','1','0','1','1','1','1','0'),
            ('0','0','0','1','0','0','1','1','1','0','0','0','0','0'),
            ('0','0','0','1','0','0','1','1','1','0','0','0','1','0'),
            ('0','0','0','1','0','0','1','1','1','0','0','1','0','0'),
            ('0','0','0','1','0','0','1','1','1','0','0','1','1','0'),
            ('0','0','0','1','0','0','1','1','1','0','1','0','0','0'),
            ('0','0','0','1','0','0','1','1','1','0','1','0','1','0'),
            ('0','0','0','1','0','0','1','1','1','0','1','1','0','0'),
            ('0','0','0','1','0','0','1','1','1','0','1','1','1','0'),
            ('0','0','0','1','0','0','1','1','1','1','0','0','0','0'),
            ('0','0','0','1','0','0','1','1','1','1','0','0','1','0'),
            ('0','0','0','1','0','0','1','1','1','1','0','1','0','0'),
            ('0','0','0','1','0','0','1','1','1','1','0','1','1','0'),
            ('0','0','0','1','0','0','1','1','1','1','1','0','0','0'),
            ('0','0','0','1','0','0','1','1','1','1','1','0','1','0'),
            ('0','0','0','1','0','0','1','1','1','1','1','1','0','0'),
            ('0','0','0','1','0','0','1','1','1','1','1','1','1','0'),
            ('0','0','0','1','0','1','0','0','0','0','0','0','0','0'),
            ('0','0','0','1','0','1','0','0','0','0','0','0','1','0'),
            ('0','0','0','1','0','1','0','0','0','0','0','1','0','0'),
            ('0','0','0','1','0','1','0','0','0','0','0','1','1','0'),
            ('0','0','0','1','0','1','0','0','0','0','1','0','0','0'),
            ('0','0','0','1','0','1','0','0','0','0','1','0','1','0'),
            ('0','0','0','1','0','1','0','0','0','0','1','1','0','0'),
            ('0','0','0','1','0','1','0','0','0','0','1','1','1','0'),
            ('0','0','0','1','0','1','0','0','0','1','0','0','0','0'),
            ('0','0','0','1','0','1','0','0','0','1','0','0','1','0'),
            ('0','0','0','1','0','1','0','0','0','1','0','1','0','0'),
            ('0','0','0','1','0','1','0','0','0','1','0','1','1','0'),
            ('0','0','0','1','0','1','0','0','0','1','1','0','0','0'),
            ('0','0','0','1','0','1','0','0','0','1','1','0','1','0'),
            ('0','0','0','1','0','1','0','0','0','1','1','1','0','0'),
            ('0','0','0','1','0','1','0','0','0','1','1','1','1','0'),
            ('0','0','0','1','0','1','0','0','1','0','0','0','0','0'),
            ('0','0','0','1','0','1','0','0','1','0','0','0','1','0'),
            ('0','0','0','1','0','1','0','0','1','0','0','1','0','0'),
            ('0','0','0','1','0','1','0','0','1','0','0','1','1','0'),
            ('0','0','0','1','0','1','0','0','1','0','1','0','0','0'),
            ('0','0','0','1','0','1','0','0','1','0','1','0','1','0'),
            ('0','0','0','1','0','1','0','0','1','0','1','1','0','0'),
            ('0','0','0','1','0','1','0','0','1','0','1','1','1','0'),
            ('0','0','0','1','0','1','0','0','1','1','0','0','0','0'),
            ('0','0','0','1','0','1','0','0','1','1','0','0','1','0'),
            ('0','0','0','1','0','1','0','0','1','1','0','1','0','0'),
            ('0','0','0','1','0','1','0','0','1','1','0','1','1','0'),
            ('0','0','0','1','0','1','0','0','1','1','1','0','0','0'),
            ('0','0','0','1','0','1','0','0','1','1','1','0','1','0'),
            ('0','0','0','1','0','1','0','0','1','1','1','1','0','0'),
            ('0','0','0','1','0','1','0','0','1','1','1','1','1','0'),
            ('0','0','0','1','0','1','0','1','0','0','0','0','0','0'),
            ('0','0','0','1','0','1','0','1','0','0','0','0','1','0'),
            ('0','0','0','1','0','1','0','1','0','0','0','1','0','0'),
            ('0','0','0','1','0','1','0','1','0','0','0','1','1','0'),
            ('0','0','0','1','0','1','0','1','0','0','1','0','0','0'),
            ('0','0','0','1','0','1','0','1','0','0','1','0','1','0'),
            ('0','0','0','1','0','1','0','1','0','0','1','1','0','0'),
            ('0','0','0','1','0','1','0','1','0','0','1','1','1','0'),
            ('0','0','0','1','0','1','0','1','0','1','0','0','0','0'),
            ('0','0','0','1','0','1','0','1','0','1','0','0','1','0'),
            ('0','0','0','1','0','1','0','1','0','1','0','1','0','0'),
            ('0','0','0','1','0','1','0','1','0','1','0','1','1','0'),
            ('0','0','0','1','0','1','0','1','0','1','1','0','0','0'),
            ('0','0','0','1','0','1','0','1','0','1','1','0','1','0'),
            ('0','0','0','1','0','1','0','1','0','1','1','1','0','0'),
            ('0','0','0','1','0','1','0','1','0','1','1','1','1','0'),
            ('0','0','0','1','0','1','0','1','1','0','0','0','0','0'),
            ('0','0','0','1','0','1','0','1','1','0','0','0','1','0'),
            ('0','0','0','1','0','1','0','1','1','0','0','1','0','0'),
            ('0','0','0','1','0','1','0','1','1','0','0','1','1','0'),
            ('0','0','0','1','0','1','0','1','1','0','1','0','0','0'),
            ('0','0','0','1','0','1','0','1','1','0','1','0','1','0'),
            ('0','0','0','1','0','1','0','1','1','0','1','1','0','0'),
            ('0','0','0','1','0','1','0','1','1','0','1','1','1','0'),
            ('0','0','0','1','0','1','0','1','1','1','0','0','0','0'),
            ('0','0','0','1','0','1','0','1','1','1','0','0','1','0'),
            ('0','0','0','1','0','1','0','1','1','1','0','1','0','0'),
            ('0','0','0','1','0','1','0','1','1','1','0','1','1','0'),
            ('0','0','0','1','0','1','0','1','1','1','1','0','0','0'),
            ('0','0','0','1','0','1','0','1','1','1','1','0','1','0'),
            ('0','0','0','1','0','1','0','1','1','1','1','1','0','0'),
            ('0','0','0','1','0','1','0','1','1','1','1','1','1','0'),
            ('0','0','0','1','0','1','1','0','0','0','0','0','0','0'),
            ('0','0','0','1','0','1','1','0','0','0','0','0','1','0'),
            ('0','0','0','1','0','1','1','0','0','0','0','1','0','0'),
            ('0','0','0','1','0','1','1','0','0','0','0','1','1','0'),
            ('0','0','0','1','0','1','1','0','0','0','1','0','0','0'),
            ('0','0','0','1','0','1','1','0','0','0','1','0','1','0'),
            ('0','0','0','1','0','1','1','0','0','0','1','1','0','0'),
            ('0','0','0','1','0','1','1','0','0','0','1','1','1','0'),
            ('0','0','0','1','0','1','1','0','0','1','0','0','0','0'),
            ('0','0','0','1','0','1','1','0','0','1','0','0','1','0'),
            ('0','0','0','1','0','1','1','0','0','1','0','1','0','0'),
            ('0','0','0','1','0','1','1','0','0','1','0','1','1','0'),
            ('0','0','0','1','0','1','1','0','0','1','1','0','0','0'),
            ('0','0','0','1','0','1','1','0','0','1','1','0','1','0'),
            ('0','0','0','1','0','1','1','0','0','1','1','1','0','0'),
            ('0','0','0','1','0','1','1','0','0','1','1','1','1','0'),
            ('0','0','0','1','0','1','1','0','1','0','0','0','0','0'),
            ('0','0','0','1','0','1','1','0','1','0','0','0','1','0'),
            ('0','0','0','1','0','1','1','0','1','0','0','1','0','0'),
            ('0','0','0','1','0','1','1','0','1','0','0','1','1','0'),
            ('0','0','0','1','0','1','1','0','1','0','1','0','0','0'),
            ('0','0','0','1','0','1','1','0','1','0','1','0','1','0'),
            ('0','0','0','1','0','1','1','0','1','0','1','1','0','0'),
            ('0','0','0','1','0','1','1','0','1','0','1','1','1','0'),
            ('0','0','0','1','0','1','1','0','1','1','0','0','0','0'),
            ('0','0','0','1','0','1','1','0','1','1','0','0','1','0'),
            ('0','0','0','1','0','1','1','0','1','1','0','1','0','0'),
            ('0','0','0','1','0','1','1','0','1','1','0','1','1','0'),
            ('0','0','0','1','0','1','1','0','1','1','1','0','0','0'),
            ('0','0','0','1','0','1','1','0','1','1','1','0','1','0'),
            ('0','0','0','1','0','1','1','0','1','1','1','1','0','0'),
            ('0','0','0','1','0','1','1','0','1','1','1','1','1','0'),
            ('0','0','0','1','0','1','1','1','0','0','0','0','0','0'),
            ('0','0','0','1','0','1','1','1','0','0','0','0','1','0'),
            ('0','0','0','1','0','1','1','1','0','0','0','1','0','0'),
            ('0','0','0','1','0','1','1','1','0','0','0','1','1','0'),
            ('0','0','0','1','0','1','1','1','0','0','1','0','0','0'),
            ('0','0','0','1','0','1','1','1','0','0','1','0','1','0'),
            ('0','0','0','1','0','1','1','1','0','0','1','1','0','0'),
            ('0','0','0','1','0','1','1','1','0','0','1','1','1','0'),
            ('0','0','0','1','0','1','1','1','0','1','0','0','0','0'),
            ('0','0','0','1','0','1','1','1','0','1','0','0','1','0'),
            ('0','0','0','1','0','1','1','1','0','1','0','1','0','0'),
            ('0','0','0','1','0','1','1','1','0','1','0','1','1','0'),
            ('0','0','0','1','0','1','1','1','0','1','1','0','0','0'),
            ('0','0','0','1','0','1','1','1','0','1','1','0','1','0'),
            ('0','0','0','1','0','1','1','1','0','1','1','1','0','0'),
            ('0','0','0','1','0','1','1','1','0','1','1','1','1','0'),
            ('0','0','0','1','0','1','1','1','1','0','0','0','0','0'),
            ('0','0','0','1','0','1','1','1','1','0','0','0','1','0'),
            ('0','0','0','1','0','1','1','1','1','0','0','1','0','0'),
            ('0','0','0','1','0','1','1','1','1','0','0','1','1','0'),
            ('0','0','0','1','0','1','1','1','1','0','1','0','0','0'),
            ('0','0','0','1','0','1','1','1','1','0','1','0','1','0'),
            ('0','0','0','1','0','1','1','1','1','0','1','1','0','0'),
            ('0','0','0','1','0','1','1','1','1','0','1','1','1','0'),
            ('0','0','0','1','0','1','1','1','1','1','0','0','0','0'),
            ('0','0','0','1','0','1','1','1','1','1','0','0','1','0'),
            ('0','0','0','1','0','1','1','1','1','1','0','1','0','0'),
            ('0','0','0','1','0','1','1','1','1','1','0','1','1','0'),
            ('0','0','0','1','0','1','1','1','1','1','1','0','0','0'),
            ('0','0','0','1','0','1','1','1','1','1','1','0','1','0'),
            ('0','0','0','1','0','1','1','1','1','1','1','1','0','0'),
            ('0','0','0','1','0','1','1','1','1','1','1','1','1','0'),
            ('0','0','0','1','1','0','0','0','0','0','0','0','0','0'),
            ('0','0','0','1','1','0','0','0','0','0','0','0','1','0'),
            ('0','0','0','1','1','0','0','0','0','0','0','1','0','0'),
            ('0','0','0','1','1','0','0','0','0','0','0','1','1','0'),
            ('0','0','0','1','1','0','0','0','0','0','1','0','0','0'),
            ('0','0','0','1','1','0','0','0','0','0','1','0','1','0'),
            ('0','0','0','1','1','0','0','0','0','0','1','1','0','0'),
            ('0','0','0','1','1','0','0','0','0','0','1','1','1','0'),
            ('0','0','0','1','1','0','0','0','0','1','0','0','0','0'),
            ('0','0','0','1','1','0','0','0','0','1','0','0','1','0'),
            ('0','0','0','1','1','0','0','0','0','1','0','1','0','0'),
            ('0','0','0','1','1','0','0','0','0','1','0','1','1','0'),
            ('0','0','0','1','1','0','0','0','0','1','1','0','0','0'),
            ('0','0','0','1','1','0','0','0','0','1','1','0','1','0'),
            ('0','0','0','1','1','0','0','0','0','1','1','1','0','0'),
            ('0','0','0','1','1','0','0','0','0','1','1','1','1','0'),
            ('0','0','0','1','1','0','0','0','1','0','0','0','0','0'),
            ('0','0','0','1','1','0','0','0','1','0','0','0','1','0'),
            ('0','0','0','1','1','0','0','0','1','0','0','1','0','0'),
            ('0','0','0','1','1','0','0','0','1','0','0','1','1','0'),
            ('0','0','0','1','1','0','0','0','1','0','1','0','0','0'),
            ('0','0','0','1','1','0','0','0','1','0','1','0','1','0'),
            ('0','0','0','1','1','0','0','0','1','0','1','1','0','0'),
            ('0','0','0','1','1','0','0','0','1','0','1','1','1','0'),
            ('0','0','0','1','1','0','0','0','1','1','0','0','0','0'),
            ('0','0','0','1','1','0','0','0','1','1','0','0','1','0'),
            ('0','0','0','1','1','0','0','0','1','1','0','1','0','0'),
            ('0','0','0','1','1','0','0','0','1','1','0','1','1','0'),
            ('0','0','0','1','1','0','0','0','1','1','1','0','0','0'),
            ('0','0','0','1','1','0','0','0','1','1','1','0','1','0'),
            ('0','0','0','1','1','0','0','0','1','1','1','1','0','0'),
            ('0','0','0','1','1','0','0','0','1','1','1','1','1','0'),
            ('0','0','0','1','1','0','0','1','0','0','0','0','0','0'),
            ('0','0','0','1','1','0','0','1','0','0','0','0','1','0'),
            ('0','0','0','1','1','0','0','1','0','0','0','1','0','0'),
            ('0','0','0','1','1','0','0','1','0','0','0','1','1','0'),
            ('0','0','0','1','1','0','0','1','0','0','1','0','0','0'),
            ('0','0','0','1','1','0','0','1','0','0','1','0','1','0'),
            ('0','0','0','1','1','0','0','1','0','0','1','1','0','0'),
            ('0','0','0','1','1','0','0','1','0','0','1','1','1','0'),
            ('0','0','0','1','1','0','0','1','0','1','0','0','0','0'),
            ('0','0','0','1','1','0','0','1','0','1','0','0','1','0'),
            ('0','0','0','1','1','0','0','1','0','1','0','1','0','0'),
            ('0','0','0','1','1','0','0','1','0','1','0','1','1','0'),
            ('0','0','0','1','1','0','0','1','0','1','1','0','0','0'),
            ('0','0','0','1','1','0','0','1','0','1','1','0','1','0'),
            ('0','0','0','1','1','0','0','1','0','1','1','1','0','0'),
            ('0','0','0','1','1','0','0','1','0','1','1','1','1','0'),
            ('0','0','0','1','1','0','0','1','1','0','0','0','0','0'),
            ('0','0','0','1','1','0','0','1','1','0','0','0','1','0'),
            ('0','0','0','1','1','0','0','1','1','0','0','1','0','0'),
            ('0','0','0','1','1','0','0','1','1','0','0','1','1','0'),
            ('0','0','0','1','1','0','0','1','1','0','1','0','0','0'),
            ('0','0','0','1','1','0','0','1','1','0','1','0','1','0'),
            ('0','0','0','1','1','0','0','1','1','0','1','1','0','0'),
            ('0','0','0','1','1','0','0','1','1','0','1','1','1','0'),
            ('0','0','0','1','1','0','0','1','1','1','0','0','0','0'),
            ('0','0','0','1','1','0','0','1','1','1','0','0','1','0'),
            ('0','0','0','1','1','0','0','1','1','1','0','1','0','0'),
            ('0','0','0','1','1','0','0','1','1','1','0','1','1','0'),
            ('0','0','0','1','1','0','0','1','1','1','1','0','0','0'),
            ('0','0','0','1','1','0','0','1','1','1','1','0','1','0'),
            ('0','0','0','1','1','0','0','1','1','1','1','1','0','0'),
            ('0','0','0','1','1','0','0','1','1','1','1','1','1','0'),
            ('0','0','0','1','1','0','1','0','0','0','0','0','0','0'),
            ('0','0','0','1','1','0','1','0','0','0','0','0','1','0'),
            ('0','0','0','1','1','0','1','0','0','0','0','1','0','0'),
            ('0','0','0','1','1','0','1','0','0','0','0','1','1','0'),
            ('0','0','0','1','1','0','1','0','0','0','1','0','0','0'),
            ('0','0','0','1','1','0','1','0','0','0','1','0','1','0'),
            ('0','0','0','1','1','0','1','0','0','0','1','1','0','0'),
            ('0','0','0','1','1','0','1','0','0','0','1','1','1','0'),
            ('0','0','0','1','1','0','1','0','0','1','0','0','0','0'),
            ('0','0','0','1','1','0','1','0','0','1','0','0','1','0'),
            ('0','0','0','1','1','0','1','0','0','1','0','1','0','0'),
            ('0','0','0','1','1','0','1','0','0','1','0','1','1','0'),
            ('0','0','0','1','1','0','1','0','0','1','1','0','0','0'),
            ('0','0','0','1','1','0','1','0','0','1','1','0','1','0'),
            ('0','0','0','1','1','0','1','0','0','1','1','1','0','0'),
            ('0','0','0','1','1','0','1','0','0','1','1','1','1','0'),
            ('0','0','0','1','1','0','1','0','1','0','0','0','0','0'),
            ('0','0','0','1','1','0','1','0','1','0','0','0','1','0'),
            ('0','0','0','1','1','0','1','0','1','0','0','1','0','0'),
            ('0','0','0','1','1','0','1','0','1','0','0','1','1','0'),
            ('0','0','0','1','1','0','1','0','1','0','1','0','0','0'),
            ('0','0','0','1','1','0','1','0','1','0','1','0','1','0'),
            ('0','0','0','1','1','0','1','0','1','0','1','1','0','0'),
            ('0','0','0','1','1','0','1','0','1','0','1','1','1','0'),
            ('0','0','0','1','1','0','1','0','1','1','0','0','0','0'),
            ('0','0','0','1','1','0','1','0','1','1','0','0','1','0'),
            ('0','0','0','1','1','0','1','0','1','1','0','1','0','0'),
            ('0','0','0','1','1','0','1','0','1','1','0','1','1','0'),
            ('0','0','0','1','1','0','1','0','1','1','1','0','0','0'),
            ('0','0','0','1','1','0','1','0','1','1','1','0','1','0'),
            ('0','0','0','1','1','0','1','0','1','1','1','1','0','0'),
            ('0','0','0','1','1','0','1','0','1','1','1','1','1','0'),
            ('0','0','0','1','1','0','1','1','0','0','0','0','0','0'),
            ('0','0','0','1','1','0','1','1','0','0','0','0','1','0'),
            ('0','0','0','1','1','0','1','1','0','0','0','1','0','0'),
            ('0','0','0','1','1','0','1','1','0','0','0','1','1','0'),
            ('0','0','0','1','1','0','1','1','0','0','1','0','0','0'),
            ('0','0','0','1','1','0','1','1','0','0','1','0','1','0'),
            ('0','0','0','1','1','0','1','1','0','0','1','1','0','0'),
            ('0','0','0','1','1','0','1','1','0','0','1','1','1','0'),
            ('0','0','0','1','1','0','1','1','0','1','0','0','0','0'),
            ('0','0','0','1','1','0','1','1','0','1','0','0','1','0'),
            ('0','0','0','1','1','0','1','1','0','1','0','1','0','0'),
            ('0','0','0','1','1','0','1','1','0','1','0','1','1','0'),
            ('0','0','0','1','1','0','1','1','0','1','1','0','0','0'),
            ('0','0','0','1','1','0','1','1','0','1','1','0','1','0'),
            ('0','0','0','1','1','0','1','1','0','1','1','1','0','0'),
            ('0','0','0','1','1','0','1','1','0','1','1','1','1','0'),
            ('0','0','0','1','1','0','1','1','1','0','0','0','0','0'),
            ('0','0','0','1','1','0','1','1','1','0','0','0','1','0'),
            ('0','0','0','1','1','0','1','1','1','0','0','1','0','0'),
            ('0','0','0','1','1','0','1','1','1','0','0','1','1','0'),
            ('0','0','0','1','1','0','1','1','1','0','1','0','0','0'),
            ('0','0','0','1','1','0','1','1','1','0','1','0','1','0'),
            ('0','0','0','1','1','0','1','1','1','0','1','1','0','0'),
            ('0','0','0','1','1','0','1','1','1','0','1','1','1','0'),
            ('0','0','0','1','1','0','1','1','1','1','0','0','0','0'),
            ('0','0','0','1','1','0','1','1','1','1','0','0','1','0'),
            ('0','0','0','1','1','0','1','1','1','1','0','1','0','0'),
            ('0','0','0','1','1','0','1','1','1','1','0','1','1','0'),
            ('0','0','0','1','1','0','1','1','1','1','1','0','0','0'),
            ('0','0','0','1','1','0','1','1','1','1','1','0','1','0'),
            ('0','0','0','1','1','0','1','1','1','1','1','1','0','0'),
            ('0','0','0','1','1','0','1','1','1','1','1','1','1','0'),
            ('0','0','0','1','1','1','0','0','0','0','0','0','0','0'),
            ('0','0','0','1','1','1','0','0','0','0','0','0','1','0'),
            ('0','0','0','1','1','1','0','0','0','0','0','1','0','0'),
            ('0','0','0','1','1','1','0','0','0','0','0','1','1','0'),
            ('0','0','0','1','1','1','0','0','0','0','1','0','0','0'),
            ('0','0','0','1','1','1','0','0','0','0','1','0','1','0'),
            ('0','0','0','1','1','1','0','0','0','0','1','1','0','0'),
            ('0','0','0','1','1','1','0','0','0','0','1','1','1','0'),
            ('0','0','0','1','1','1','0','0','0','1','0','0','0','0'),
            ('0','0','0','1','1','1','0','0','0','1','0','0','1','0'),
            ('0','0','0','1','1','1','0','0','0','1','0','1','0','0'),
            ('0','0','0','1','1','1','0','0','0','1','0','1','1','0'),
            ('0','0','0','1','1','1','0','0','0','1','1','0','0','0'),
            ('0','0','0','1','1','1','0','0','0','1','1','0','1','0'),
            ('0','0','0','1','1','1','0','0','0','1','1','1','0','0'),
            ('0','0','0','1','1','1','0','0','0','1','1','1','1','0'),
            ('0','0','0','1','1','1','0','0','1','0','0','0','0','0'),
            ('0','0','0','1','1','1','0','0','1','0','0','0','1','0'),
            ('0','0','0','1','1','1','0','0','1','0','0','1','0','0'),
            ('0','0','0','1','1','1','0','0','1','0','0','1','1','0'),
            ('0','0','0','1','1','1','0','0','1','0','1','0','0','0'),
            ('0','0','0','1','1','1','0','0','1','0','1','0','1','0'),
            ('0','0','0','1','1','1','0','0','1','0','1','1','0','0'),
            ('0','0','0','1','1','1','0','0','1','0','1','1','1','0'),
            ('0','0','0','1','1','1','0','0','1','1','0','0','0','0'),
            ('0','0','0','1','1','1','0','0','1','1','0','0','1','0'),
            ('0','0','0','1','1','1','0','0','1','1','0','1','0','0'),
            ('0','0','0','1','1','1','0','0','1','1','0','1','1','0'),
            ('0','0','0','1','1','1','0','0','1','1','1','0','0','0'),
            ('0','0','0','1','1','1','0','0','1','1','1','0','1','0'),
            ('0','0','0','1','1','1','0','0','1','1','1','1','0','0'),
            ('0','0','0','1','1','1','0','0','1','1','1','1','1','0'),
            ('0','0','0','1','1','1','0','1','0','0','0','0','0','0'),
            ('0','0','0','1','1','1','0','1','0','0','0','0','1','0'),
            ('0','0','0','1','1','1','0','1','0','0','0','1','0','0'),
            ('0','0','0','1','1','1','0','1','0','0','0','1','1','0'),
            ('0','0','0','1','1','1','0','1','0','0','1','0','0','0'),
            ('0','0','0','1','1','1','0','1','0','0','1','0','1','0'),
            ('0','0','0','1','1','1','0','1','0','0','1','1','0','0'),
            ('0','0','0','1','1','1','0','1','0','0','1','1','1','0'),
            ('0','0','0','1','1','1','0','1','0','1','0','0','0','0'),
            ('0','0','0','1','1','1','0','1','0','1','0','0','1','0'),
            ('0','0','0','1','1','1','0','1','0','1','0','1','0','0'),
            ('0','0','0','1','1','1','0','1','0','1','0','1','1','0'),
            ('0','0','0','1','1','1','0','1','0','1','1','0','0','0'),
            ('0','0','0','1','1','1','0','1','0','1','1','0','1','0'),
            ('0','0','0','1','1','1','0','1','0','1','1','1','0','0'),
            ('0','0','0','1','1','1','0','1','0','1','1','1','1','0'),
            ('0','0','0','1','1','1','0','1','1','0','0','0','0','0'),
            ('0','0','0','1','1','1','0','1','1','0','0','0','1','0'),
            ('0','0','0','1','1','1','0','1','1','0','0','1','0','0'),
            ('0','0','0','1','1','1','0','1','1','0','0','1','1','0'),
            ('0','0','0','1','1','1','0','1','1','0','1','0','0','0'),
            ('0','0','0','1','1','1','0','1','1','0','1','0','1','0'),
            ('0','0','0','1','1','1','0','1','1','0','1','1','0','0'),
            ('0','0','0','1','1','1','0','1','1','0','1','1','1','0'),
            ('0','0','0','1','1','1','0','1','1','1','0','0','0','0'),
            ('0','0','0','1','1','1','0','1','1','1','0','0','1','0'),
            ('0','0','0','1','1','1','0','1','1','1','0','1','0','0'),
            ('0','0','0','1','1','1','0','1','1','1','0','1','1','0'),
            ('0','0','0','1','1','1','0','1','1','1','1','0','0','0'),
            ('0','0','0','1','1','1','0','1','1','1','1','0','1','0'),
            ('0','0','0','1','1','1','0','1','1','1','1','1','0','0'),
            ('0','0','0','1','1','1','0','1','1','1','1','1','1','0'),
            ('0','0','0','1','1','1','1','0','0','0','0','0','0','0'),
            ('0','0','0','1','1','1','1','0','0','0','0','0','1','0'),
            ('0','0','0','1','1','1','1','0','0','0','0','1','0','0'),
            ('0','0','0','1','1','1','1','0','0','0','0','1','1','0'),
            ('0','0','0','1','1','1','1','0','0','0','1','0','0','0'),
            ('0','0','0','1','1','1','1','0','0','0','1','0','1','0'),
            ('0','0','0','1','1','1','1','0','0','0','1','1','0','0'),
            ('0','0','0','1','1','1','1','0','0','0','1','1','1','0'),
            ('0','0','0','1','1','1','1','0','0','1','0','0','0','0'),
            ('0','0','0','1','1','1','1','0','0','1','0','0','1','0'),
            ('0','0','0','1','1','1','1','0','0','1','0','1','0','0'),
            ('0','0','0','1','1','1','1','0','0','1','0','1','1','0'),
            ('0','0','0','1','1','1','1','0','0','1','1','0','0','0'),
            ('0','0','0','1','1','1','1','0','0','1','1','0','1','0'),
            ('0','0','0','1','1','1','1','0','0','1','1','1','0','0'),
            ('0','0','0','1','1','1','1','0','0','1','1','1','1','0'),
            ('0','0','0','1','1','1','1','0','1','0','0','0','0','0'),
            ('0','0','0','1','1','1','1','0','1','0','0','0','1','0'),
            ('0','0','0','1','1','1','1','0','1','0','0','1','0','0'),
            ('0','0','0','1','1','1','1','0','1','0','0','1','1','0'),
            ('0','0','0','1','1','1','1','0','1','0','1','0','0','0'),
            ('0','0','0','1','1','1','1','0','1','0','1','0','1','0'),
            ('0','0','0','1','1','1','1','0','1','0','1','1','0','0'),
            ('0','0','0','1','1','1','1','0','1','0','1','1','1','0'),
            ('0','0','0','1','1','1','1','0','1','1','0','0','0','0'),
            ('0','0','0','1','1','1','1','0','1','1','0','0','1','0'),
            ('0','0','0','1','1','1','1','0','1','1','0','1','0','0'),
            ('0','0','0','1','1','1','1','0','1','1','0','1','1','0'),
            ('0','0','0','1','1','1','1','0','1','1','1','0','0','0'),
            ('0','0','0','1','1','1','1','0','1','1','1','0','1','0'),
            ('0','0','0','1','1','1','1','0','1','1','1','1','0','0'),
            ('0','0','0','1','1','1','1','0','1','1','1','1','1','0'),
            ('0','0','0','1','1','1','1','1','0','0','0','0','0','0'),
            ('0','0','0','1','1','1','1','1','0','0','0','0','1','0'),
            ('0','0','0','1','1','1','1','1','0','0','0','1','0','0'),
            ('0','0','0','1','1','1','1','1','0','0','0','1','1','0'),
            ('0','0','0','1','1','1','1','1','0','0','1','0','0','0'),
            ('0','0','0','1','1','1','1','1','0','0','1','0','1','0'),
            ('0','0','0','1','1','1','1','1','0','0','1','1','0','0'),
            ('0','0','0','1','1','1','1','1','0','0','1','1','1','0'),
            ('0','0','0','1','1','1','1','1','0','1','0','0','0','0'),
            ('0','0','0','1','1','1','1','1','0','1','0','0','1','0'),
            ('0','0','0','1','1','1','1','1','0','1','0','1','0','0'),
            ('0','0','0','1','1','1','1','1','0','1','0','1','1','0'),
            ('0','0','0','1','1','1','1','1','0','1','1','0','0','0'),
            ('0','0','0','1','1','1','1','1','0','1','1','0','1','0'),
            ('0','0','0','1','1','1','1','1','0','1','1','1','0','0'),
            ('0','0','0','1','1','1','1','1','0','1','1','1','1','0'),
            ('0','0','0','1','1','1','1','1','1','0','0','0','0','0'),
            ('0','0','0','1','1','1','1','1','1','0','0','0','1','0'),
            ('0','0','0','1','1','1','1','1','1','0','0','1','0','0'),
            ('0','0','0','1','1','1','1','1','1','0','0','1','1','0'),
            ('0','0','0','1','1','1','1','1','1','0','1','0','0','0'),
            ('0','0','0','1','1','1','1','1','1','0','1','0','1','0'),
            ('0','0','0','1','1','1','1','1','1','0','1','1','0','0'),
            ('0','0','0','1','1','1','1','1','1','0','1','1','1','0'),
            ('0','0','0','1','1','1','1','1','1','1','0','0','0','0'),
            ('0','0','0','1','1','1','1','1','1','1','0','0','1','0'),
            ('0','0','0','1','1','1','1','1','1','1','0','1','0','0'),
            ('0','0','0','1','1','1','1','1','1','1','0','1','1','0'),
            ('0','0','0','1','1','1','1','1','1','1','1','0','0','0'),
            ('0','0','0','1','1','1','1','1','1','1','1','0','1','0'),
            ('0','0','0','1','1','1','1','1','1','1','1','1','0','0'),
            ('0','0','0','1','1','1','1','1','1','1','1','1','1','0'),
            ('0','0','1','0','0','0','0','0','0','0','0','0','0','0'),
            ('0','0','1','0','0','0','0','0','0','0','0','0','1','0'),
            ('0','0','1','0','0','0','0','0','0','0','0','1','0','0'),
            ('0','0','1','0','0','0','0','0','0','0','0','1','1','0'),
            ('0','0','1','0','0','0','0','0','0','0','1','0','0','0'),
            ('0','0','1','0','0','0','0','0','0','0','1','0','1','0'),
            ('0','0','1','0','0','0','0','0','0','0','1','1','0','0'),
            ('0','0','1','0','0','0','0','0','0','0','1','1','1','0'),
            ('0','0','1','0','0','0','0','0','0','1','0','0','0','0'),
            ('0','0','1','0','0','0','0','0','0','1','0','0','1','0'),
            ('0','0','1','0','0','0','0','0','0','1','0','1','0','0'),
            ('0','0','1','0','0','0','0','0','0','1','0','1','1','0'),
            ('0','0','1','0','0','0','0','0','0','1','1','0','0','0'),
            ('0','0','1','0','0','0','0','0','0','1','1','0','1','0'),
            ('0','0','1','0','0','0','0','0','0','1','1','1','0','0'),
            ('0','0','1','0','0','0','0','0','0','1','1','1','1','0'),
            ('0','0','1','0','0','0','0','0','1','0','0','0','0','0'),
            ('0','0','1','0','0','0','0','0','1','0','0','0','1','0'),
            ('0','0','1','0','0','0','0','0','1','0','0','1','0','0'),
            ('0','0','1','0','0','0','0','0','1','0','0','1','1','0'),
            ('0','0','1','0','0','0','0','0','1','0','1','0','0','0'),
            ('0','0','1','0','0','0','0','0','1','0','1','0','1','0'),
            ('0','0','1','0','0','0','0','0','1','0','1','1','0','0'),
            ('0','0','1','0','0','0','0','0','1','0','1','1','1','0'),
            ('0','0','1','0','0','0','0','0','1','1','0','0','0','0'),
            ('0','0','1','0','0','0','0','0','1','1','0','0','1','0'),
            ('0','0','1','0','0','0','0','0','1','1','0','1','0','0'),
            ('0','0','1','0','0','0','0','0','1','1','0','1','1','0'),
            ('0','0','1','0','0','0','0','0','1','1','1','0','0','0'),
            ('0','0','1','0','0','0','0','0','1','1','1','0','1','0'),
            ('0','0','1','0','0','0','0','0','1','1','1','1','0','0'),
            ('0','0','1','0','0','0','0','0','1','1','1','1','1','0'),
            ('0','0','1','0','0','0','0','1','0','0','0','0','0','0'),
            ('0','0','1','0','0','0','0','1','0','0','0','0','1','0'),
            ('0','0','1','0','0','0','0','1','0','0','0','1','0','0'),
            ('0','0','1','0','0','0','0','1','0','0','0','1','1','0'),
            ('0','0','1','0','0','0','0','1','0','0','1','0','0','0'),
            ('0','0','1','0','0','0','0','1','0','0','1','0','1','0'),
            ('0','0','1','0','0','0','0','1','0','0','1','1','0','0'),
            ('0','0','1','0','0','0','0','1','0','0','1','1','1','0'),
            ('0','0','1','0','0','0','0','1','0','1','0','0','0','0'),
            ('0','0','1','0','0','0','0','1','0','1','0','0','1','0'),
            ('0','0','1','0','0','0','0','1','0','1','0','1','0','0'),
            ('0','0','1','0','0','0','0','1','0','1','0','1','1','0'),
            ('0','0','1','0','0','0','0','1','0','1','1','0','0','0'),
            ('0','0','1','0','0','0','0','1','0','1','1','0','1','0'),
            ('0','0','1','0','0','0','0','1','0','1','1','1','0','0'),
            ('0','0','1','0','0','0','0','1','0','1','1','1','1','0'),
            ('0','0','1','0','0','0','0','1','1','0','0','0','0','0'),
            ('0','0','1','0','0','0','0','1','1','0','0','0','1','0'),
            ('0','0','1','0','0','0','0','1','1','0','0','1','0','0'),
            ('0','0','1','0','0','0','0','1','1','0','0','1','1','0'),
            ('0','0','1','0','0','0','0','1','1','0','1','0','0','0'),
            ('0','0','1','0','0','0','0','1','1','0','1','0','1','0'),
            ('0','0','1','0','0','0','0','1','1','0','1','1','0','0'),
            ('0','0','1','0','0','0','0','1','1','0','1','1','1','0'),
            ('0','0','1','0','0','0','0','1','1','1','0','0','0','0'),
            ('0','0','1','0','0','0','0','1','1','1','0','0','1','0'),
            ('0','0','1','0','0','0','0','1','1','1','0','1','0','0'),
            ('0','0','1','0','0','0','0','1','1','1','0','1','1','0'),
            ('0','0','1','0','0','0','0','1','1','1','1','0','0','0'),
            ('0','0','1','0','0','0','0','1','1','1','1','0','1','0'),
            ('0','0','1','0','0','0','0','1','1','1','1','1','0','0'),
            ('0','0','1','0','0','0','0','1','1','1','1','1','1','0'),
            ('0','0','1','0','0','0','1','0','0','0','0','0','0','0'),
            ('0','0','1','0','0','0','1','0','0','0','0','0','1','0'),
            ('0','0','1','0','0','0','1','0','0','0','0','1','0','0'),
            ('0','0','1','0','0','0','1','0','0','0','0','1','1','0'),
            ('0','0','1','0','0','0','1','0','0','0','1','0','0','0'),
            ('0','0','1','0','0','0','1','0','0','0','1','0','1','0'),
            ('0','0','1','0','0','0','1','0','0','0','1','1','0','0'),
            ('0','0','1','0','0','0','1','0','0','0','1','1','1','0'),
            ('0','0','1','0','0','0','1','0','0','1','0','0','0','0'),
            ('0','0','1','0','0','0','1','0','0','1','0','0','1','0'),
            ('0','0','1','0','0','0','1','0','0','1','0','1','0','0'),
            ('0','0','1','0','0','0','1','0','0','1','0','1','1','0'),
            ('0','0','1','0','0','0','1','0','0','1','1','0','0','0'),
            ('0','0','1','0','0','0','1','0','0','1','1','0','1','0'),
            ('0','0','1','0','0','0','1','0','0','1','1','1','0','0'),
            ('0','0','1','0','0','0','1','0','0','1','1','1','1','0'),
            ('0','0','1','0','0','0','1','0','1','0','0','0','0','0'),
            ('0','0','1','0','0','0','1','0','1','0','0','0','1','0'),
            ('0','0','1','0','0','0','1','0','1','0','0','1','0','0'),
            ('0','0','1','0','0','0','1','0','1','0','0','1','1','0'),
            ('0','0','1','0','0','0','1','0','1','0','1','0','0','0'),
            ('0','0','1','0','0','0','1','0','1','0','1','0','1','0'),
            ('0','0','1','0','0','0','1','0','1','0','1','1','0','0'),
            ('0','0','1','0','0','0','1','0','1','0','1','1','1','0'),
            ('0','0','1','0','0','0','1','0','1','1','0','0','0','0'),
            ('0','0','1','0','0','0','1','0','1','1','0','0','1','0'),
            ('0','0','1','0','0','0','1','0','1','1','0','1','0','0'),
            ('0','0','1','0','0','0','1','0','1','1','0','1','1','0'),
            ('0','0','1','0','0','0','1','0','1','1','1','0','0','0'),
            ('0','0','1','0','0','0','1','0','1','1','1','0','1','0'),
            ('0','0','1','0','0','0','1','0','1','1','1','1','0','0'),
            ('0','0','1','0','0','0','1','0','1','1','1','1','1','0'),
            ('0','0','1','0','0','0','1','1','0','0','0','0','0','0'),
            ('0','0','1','0','0','0','1','1','0','0','0','0','1','0'),
            ('0','0','1','0','0','0','1','1','0','0','0','1','0','0'),
            ('0','0','1','0','0','0','1','1','0','0','0','1','1','0'),
            ('0','0','1','0','0','0','1','1','0','0','1','0','0','0'),
            ('0','0','1','0','0','0','1','1','0','0','1','0','1','0'),
            ('0','0','1','0','0','0','1','1','0','0','1','1','0','0'),
            ('0','0','1','0','0','0','1','1','0','0','1','1','1','0'),
            ('0','0','1','0','0','0','1','1','0','1','0','0','0','0'),
            ('0','0','1','0','0','0','1','1','0','1','0','0','1','0'),
            ('0','0','1','0','0','0','1','1','0','1','0','1','0','0'),
            ('0','0','1','0','0','0','1','1','0','1','0','1','1','0'),
            ('0','0','1','0','0','0','1','1','0','1','1','0','0','0'),
            ('0','0','1','0','0','0','1','1','0','1','1','0','1','0'),
            ('0','0','1','0','0','0','1','1','0','1','1','1','0','0'),
            ('0','0','1','0','0','0','1','1','0','1','1','1','1','0'),
            ('0','0','1','0','0','0','1','1','1','0','0','0','0','0'),
            ('0','0','1','0','0','0','1','1','1','0','0','0','1','0'),
            ('0','0','1','0','0','0','1','1','1','0','0','1','0','0'),
            ('0','0','1','0','0','0','1','1','1','0','0','1','1','0'),
            ('0','0','1','0','0','0','1','1','1','0','1','0','0','0'),
            ('0','0','1','0','0','0','1','1','1','0','1','0','1','0'),
            ('0','0','1','0','0','0','1','1','1','0','1','1','0','0'),
            ('0','0','1','0','0','0','1','1','1','0','1','1','1','0'),
            ('0','0','1','0','0','0','1','1','1','1','0','0','0','0'),
            ('0','0','1','0','0','0','1','1','1','1','0','0','1','0'),
            ('0','0','1','0','0','0','1','1','1','1','0','1','0','0'),
            ('0','0','1','0','0','0','1','1','1','1','0','1','1','0'),
            ('0','0','1','0','0','0','1','1','1','1','1','0','0','0'),
            ('0','0','1','0','0','0','1','1','1','1','1','0','1','0'),
            ('0','0','1','0','0','0','1','1','1','1','1','1','0','0'),
            ('0','0','1','0','0','0','1','1','1','1','1','1','1','0'),
            ('0','0','1','0','0','1','0','0','0','0','0','0','0','0'),
            ('0','0','1','0','0','1','0','0','0','0','0','0','1','0'),
            ('0','0','1','0','0','1','0','0','0','0','0','1','0','0'),
            ('0','0','1','0','0','1','0','0','0','0','0','1','1','0'),
            ('0','0','1','0','0','1','0','0','0','0','1','0','0','0'),
            ('0','0','1','0','0','1','0','0','0','0','1','0','1','0'),
            ('0','0','1','0','0','1','0','0','0','0','1','1','0','0'),
            ('0','0','1','0','0','1','0','0','0','0','1','1','1','0'),
            ('0','0','1','0','0','1','0','0','0','1','0','0','0','0'),
            ('0','0','1','0','0','1','0','0','0','1','0','0','1','0'),
            ('0','0','1','0','0','1','0','0','0','1','0','1','0','0'),
            ('0','0','1','0','0','1','0','0','0','1','0','1','1','0'),
            ('0','0','1','0','0','1','0','0','0','1','1','0','0','0'),
            ('0','0','1','0','0','1','0','0','0','1','1','0','1','0'),
            ('0','0','1','0','0','1','0','0','0','1','1','1','0','0'),
            ('0','0','1','0','0','1','0','0','0','1','1','1','1','0'),
            ('0','0','1','0','0','1','0','0','1','0','0','0','0','0'),
            ('0','0','1','0','0','1','0','0','1','0','0','0','1','0'),
            ('0','0','1','0','0','1','0','0','1','0','0','1','0','0'),
            ('0','0','1','0','0','1','0','0','1','0','0','1','1','0'),
            ('0','0','1','0','0','1','0','0','1','0','1','0','0','0'),
            ('0','0','1','0','0','1','0','0','1','0','1','0','1','0'),
            ('0','0','1','0','0','1','0','0','1','0','1','1','0','0'),
            ('0','0','1','0','0','1','0','0','1','0','1','1','1','0'),
            ('0','0','1','0','0','1','0','0','1','1','0','0','0','0'),
            ('0','0','1','0','0','1','0','0','1','1','0','0','1','0'),
            ('0','0','1','0','0','1','0','0','1','1','0','1','0','0'),
            ('0','0','1','0','0','1','0','0','1','1','0','1','1','0'),
            ('0','0','1','0','0','1','0','0','1','1','1','0','0','0'),
            ('0','0','1','0','0','1','0','0','1','1','1','0','1','0'),
            ('0','0','1','0','0','1','0','0','1','1','1','1','0','0'),
            ('0','0','1','0','0','1','0','0','1','1','1','1','1','0'),
            ('0','0','1','0','0','1','0','1','0','0','0','0','0','0'),
            ('0','0','1','0','0','1','0','1','0','0','0','0','1','0'),
            ('0','0','1','0','0','1','0','1','0','0','0','1','0','0'),
            ('0','0','1','0','0','1','0','1','0','0','0','1','1','0'),
            ('0','0','1','0','0','1','0','1','0','0','1','0','0','0'),
            ('0','0','1','0','0','1','0','1','0','0','1','0','1','0'),
            ('0','0','1','0','0','1','0','1','0','0','1','1','0','0'),
            ('0','0','1','0','0','1','0','1','0','0','1','1','1','0'),
            ('0','0','1','0','0','1','0','1','0','1','0','0','0','0'),
            ('0','0','1','0','0','1','0','1','0','1','0','0','1','0'),
            ('0','0','1','0','0','1','0','1','0','1','0','1','0','0'),
            ('0','0','1','0','0','1','0','1','0','1','0','1','1','0'),
            ('0','0','1','0','0','1','0','1','0','1','1','0','0','0'),
            ('0','0','1','0','0','1','0','1','0','1','1','0','1','0'),
            ('0','0','1','0','0','1','0','1','0','1','1','1','0','0'),
            ('0','0','1','0','0','1','0','1','0','1','1','1','1','0'),
            ('0','0','1','0','0','1','0','1','1','0','0','0','0','0'),
            ('0','0','1','0','0','1','0','1','1','0','0','0','1','0'),
            ('0','0','1','0','0','1','0','1','1','0','0','1','0','0'),
            ('0','0','1','0','0','1','0','1','1','0','0','1','1','0'),
            ('0','0','1','0','0','1','0','1','1','0','1','0','0','0'),
            ('0','0','1','0','0','1','0','1','1','0','1','0','1','0'),
            ('0','0','1','0','0','1','0','1','1','0','1','1','0','0'),
            ('0','0','1','0','0','1','0','1','1','0','1','1','1','0'),
            ('0','0','1','0','0','1','0','1','1','1','0','0','0','0'),
            ('0','0','1','0','0','1','0','1','1','1','0','0','1','0'),
            ('0','0','1','0','0','1','0','1','1','1','0','1','0','0'),
            ('0','0','1','0','0','1','0','1','1','1','0','1','1','0'),
            ('0','0','1','0','0','1','0','1','1','1','1','0','0','0'),
            ('0','0','1','0','0','1','0','1','1','1','1','0','1','0'),
            ('0','0','1','0','0','1','0','1','1','1','1','1','0','0'),
            ('0','0','1','0','0','1','0','1','1','1','1','1','1','0'),
            ('0','0','1','0','0','1','1','0','0','0','0','0','0','0'),
            ('0','0','1','0','0','1','1','0','0','0','0','0','1','0'),
            ('0','0','1','0','0','1','1','0','0','0','0','1','0','0'),
            ('0','0','1','0','0','1','1','0','0','0','0','1','1','0'),
            ('0','0','1','0','0','1','1','0','0','0','1','0','0','0'),
            ('0','0','1','0','0','1','1','0','0','0','1','0','1','0'),
            ('0','0','1','0','0','1','1','0','0','0','1','1','0','0'),
            ('0','0','1','0','0','1','1','0','0','0','1','1','1','0'),
            ('0','0','1','0','0','1','1','0','0','1','0','0','0','0'),
            ('0','0','1','0','0','1','1','0','0','1','0','0','1','0'),
            ('0','0','1','0','0','1','1','0','0','1','0','1','0','0'),
            ('0','0','1','0','0','1','1','0','0','1','0','1','1','0'),
            ('0','0','1','0','0','1','1','0','0','1','1','0','0','0'),
            ('0','0','1','0','0','1','1','0','0','1','1','0','1','0'),
            ('0','0','1','0','0','1','1','0','0','1','1','1','0','0'),
            ('0','0','1','0','0','1','1','0','0','1','1','1','1','0'),
            ('0','0','1','0','0','1','1','0','1','0','0','0','0','0'),
            ('0','0','1','0','0','1','1','0','1','0','0','0','1','0'),
            ('0','0','1','0','0','1','1','0','1','0','0','1','0','0'),
            ('0','0','1','0','0','1','1','0','1','0','0','1','1','0'),
            ('0','0','1','0','0','1','1','0','1','0','1','0','0','0'),
            ('0','0','1','0','0','1','1','0','1','0','1','0','1','0'),
            ('0','0','1','0','0','1','1','0','1','0','1','1','0','0'),
            ('0','0','1','0','0','1','1','0','1','0','1','1','1','0'),
            ('0','0','1','0','0','1','1','0','1','1','0','0','0','0'),
            ('0','0','1','0','0','1','1','0','1','1','0','0','1','0'),
            ('0','0','1','0','0','1','1','0','1','1','0','1','0','0'),
            ('0','0','1','0','0','1','1','0','1','1','0','1','1','0'),
            ('0','0','1','0','0','1','1','0','1','1','1','0','0','0'),
            ('0','0','1','0','0','1','1','0','1','1','1','0','1','0'),
            ('0','0','1','0','0','1','1','0','1','1','1','1','0','0'),
            ('0','0','1','0','0','1','1','0','1','1','1','1','1','0'),
            ('0','0','1','0','0','1','1','1','0','0','0','0','0','0'),
            ('0','0','1','0','0','1','1','1','0','0','0','0','1','0'),
            ('0','0','1','0','0','1','1','1','0','0','0','1','0','0'),
            ('0','0','1','0','0','1','1','1','0','0','0','1','1','0'),
            ('0','0','1','0','0','1','1','1','0','0','1','0','0','0'),
            ('0','0','1','0','0','1','1','1','0','0','1','0','1','0'),
            ('0','0','1','0','0','1','1','1','0','0','1','1','0','0'),
            ('0','0','1','0','0','1','1','1','0','0','1','1','1','0'),
            ('0','0','1','0','0','1','1','1','0','1','0','0','0','0'),
            ('0','0','1','0','0','1','1','1','0','1','0','0','1','0'),
            ('0','0','1','0','0','1','1','1','0','1','0','1','0','0'),
            ('0','0','1','0','0','1','1','1','0','1','0','1','1','0'),
            ('0','0','1','0','0','1','1','1','0','1','1','0','0','0'),
            ('0','0','1','0','0','1','1','1','0','1','1','0','1','0'),
            ('0','0','1','0','0','1','1','1','0','1','1','1','0','0'),
            ('0','0','1','0','0','1','1','1','0','1','1','1','1','0'),
            ('0','0','1','0','0','1','1','1','1','0','0','0','0','0'),
            ('0','0','1','0','0','1','1','1','1','0','0','0','1','0'),
            ('0','0','1','0','0','1','1','1','1','0','0','1','0','0'),
            ('0','0','1','0','0','1','1','1','1','0','0','1','1','0'),
            ('0','0','1','0','0','1','1','1','1','0','1','0','0','0'),
            ('0','0','1','0','0','1','1','1','1','0','1','0','1','0'),
            ('0','0','1','0','0','1','1','1','1','0','1','1','0','0'),
            ('0','0','1','0','0','1','1','1','1','0','1','1','1','0'),
            ('0','0','1','0','0','1','1','1','1','1','0','0','0','0'),
            ('0','0','1','0','0','1','1','1','1','1','0','0','1','0'),
            ('0','0','1','0','0','1','1','1','1','1','0','1','0','0'),
            ('0','0','1','0','0','1','1','1','1','1','0','1','1','0'),
            ('0','0','1','0','0','1','1','1','1','1','1','0','0','0'),
            ('0','0','1','0','0','1','1','1','1','1','1','0','1','0'),
            ('0','0','1','0','0','1','1','1','1','1','1','1','0','0'),
            ('0','0','1','0','0','1','1','1','1','1','1','1','1','0'),
            ('0','0','1','0','1','0','0','0','0','0','0','0','0','0'),
            ('0','0','1','0','1','0','0','0','0','0','0','0','1','0'),
            ('0','0','1','0','1','0','0','0','0','0','0','1','0','0'),
            ('0','0','1','0','1','0','0','0','0','0','0','1','1','0'),
            ('0','0','1','0','1','0','0','0','0','0','1','0','0','0'),
            ('0','0','1','0','1','0','0','0','0','0','1','0','1','0'),
            ('0','0','1','0','1','0','0','0','0','0','1','1','0','0'),
            ('0','0','1','0','1','0','0','0','0','0','1','1','1','0'),
            ('0','0','1','0','1','0','0','0','0','1','0','0','0','0'),
            ('0','0','1','0','1','0','0','0','0','1','0','0','1','0'),
            ('0','0','1','0','1','0','0','0','0','1','0','1','0','0'),
            ('0','0','1','0','1','0','0','0','0','1','0','1','1','0'),
            ('0','0','1','0','1','0','0','0','0','1','1','0','0','0'),
            ('0','0','1','0','1','0','0','0','0','1','1','0','1','0'),
            ('0','0','1','0','1','0','0','0','0','1','1','1','0','0'),
            ('0','0','1','0','1','0','0','0','0','1','1','1','1','0'),
            ('0','0','1','0','1','0','0','0','1','0','0','0','0','0'),
            ('0','0','1','0','1','0','0','0','1','0','0','0','1','0'),
            ('0','0','1','0','1','0','0','0','1','0','0','1','0','0'),
            ('0','0','1','0','1','0','0','0','1','0','0','1','1','0'),
            ('0','0','1','0','1','0','0','0','1','0','1','0','0','0'),
            ('0','0','1','0','1','0','0','0','1','0','1','0','1','0'),
            ('0','0','1','0','1','0','0','0','1','0','1','1','0','0'),
            ('0','0','1','0','1','0','0','0','1','0','1','1','1','0'),
            ('0','0','1','0','1','0','0','0','1','1','0','0','0','0'),
            ('0','0','1','0','1','0','0','0','1','1','0','0','1','0'),
            ('0','0','1','0','1','0','0','0','1','1','0','1','0','0'),
            ('0','0','1','0','1','0','0','0','1','1','0','1','1','0'),
            ('0','0','1','0','1','0','0','0','1','1','1','0','0','0'),
            ('0','0','1','0','1','0','0','0','1','1','1','0','1','0'),
            ('0','0','1','0','1','0','0','0','1','1','1','1','0','0'),
            ('0','0','1','0','1','0','0','0','1','1','1','1','1','0'),
            ('0','0','1','0','1','0','0','1','0','0','0','0','0','0'),
            ('0','0','1','0','1','0','0','1','0','0','0','0','1','0'),
            ('0','0','1','0','1','0','0','1','0','0','0','1','0','0'),
            ('0','0','1','0','1','0','0','1','0','0','0','1','1','0'),
            ('0','0','1','0','1','0','0','1','0','0','1','0','0','0'),
            ('0','0','1','0','1','0','0','1','0','0','1','0','1','0'),
            ('0','0','1','0','1','0','0','1','0','0','1','1','0','0'),
            ('0','0','1','0','1','0','0','1','0','0','1','1','1','0'),
            ('0','0','1','0','1','0','0','1','0','1','0','0','0','0'),
            ('0','0','1','0','1','0','0','1','0','1','0','0','1','0'),
            ('0','0','1','0','1','0','0','1','0','1','0','1','0','0'),
            ('0','0','1','0','1','0','0','1','0','1','0','1','1','0'),
            ('0','0','1','0','1','0','0','1','0','1','1','0','0','0'),
            ('0','0','1','0','1','0','0','1','0','1','1','0','1','0'),
            ('0','0','1','0','1','0','0','1','0','1','1','1','0','0'),
            ('0','0','1','0','1','0','0','1','0','1','1','1','1','0'),
            ('0','0','1','0','1','0','0','1','1','0','0','0','0','0'),
            ('0','0','1','0','1','0','0','1','1','0','0','0','1','0'),
            ('0','0','1','0','1','0','0','1','1','0','0','1','0','0'),
            ('0','0','1','0','1','0','0','1','1','0','0','1','1','0'),
            ('0','0','1','0','1','0','0','1','1','0','1','0','0','0'),
            ('0','0','1','0','1','0','0','1','1','0','1','0','1','0'),
            ('0','0','1','0','1','0','0','1','1','0','1','1','0','0'),
            ('0','0','1','0','1','0','0','1','1','0','1','1','1','0'),
            ('0','0','1','0','1','0','0','1','1','1','0','0','0','0'),
            ('0','0','1','0','1','0','0','1','1','1','0','0','1','0'),
            ('0','0','1','0','1','0','0','1','1','1','0','1','0','0'),
            ('0','0','1','0','1','0','0','1','1','1','0','1','1','0'),
            ('0','0','1','0','1','0','0','1','1','1','1','0','0','0'),
            ('0','0','1','0','1','0','0','1','1','1','1','0','1','0'),
            ('0','0','1','0','1','0','0','1','1','1','1','1','0','0'),
            ('0','0','1','0','1','0','0','1','1','1','1','1','1','0'),
            ('0','0','1','0','1','0','1','0','0','0','0','0','0','0'),
            ('0','0','1','0','1','0','1','0','0','0','0','0','1','0'),
            ('0','0','1','0','1','0','1','0','0','0','0','1','0','0'),
            ('0','0','1','0','1','0','1','0','0','0','0','1','1','0'),
            ('0','0','1','0','1','0','1','0','0','0','1','0','0','0'),
            ('0','0','1','0','1','0','1','0','0','0','1','0','1','0'),
            ('0','0','1','0','1','0','1','0','0','0','1','1','0','0'),
            ('0','0','1','0','1','0','1','0','0','0','1','1','1','0'),
            ('0','0','1','0','1','0','1','0','0','1','0','0','0','0'),
            ('0','0','1','0','1','0','1','0','0','1','0','0','1','0'),
            ('0','0','1','0','1','0','1','0','0','1','0','1','0','0'),
            ('0','0','1','0','1','0','1','0','0','1','0','1','1','0'),
            ('0','0','1','0','1','0','1','0','0','1','1','0','0','0'),
            ('0','0','1','0','1','0','1','0','0','1','1','0','1','0'),
            ('0','0','1','0','1','0','1','0','0','1','1','1','0','0'),
            ('0','0','1','0','1','0','1','0','0','1','1','1','1','0'),
            ('0','0','1','0','1','0','1','0','1','0','0','0','0','0'),
            ('0','0','1','0','1','0','1','0','1','0','0','0','1','0'),
            ('0','0','1','0','1','0','1','0','1','0','0','1','0','0'),
            ('0','0','1','0','1','0','1','0','1','0','0','1','1','0'),
            ('0','0','1','0','1','0','1','0','1','0','1','0','0','0'),
            ('0','0','1','0','1','0','1','0','1','0','1','0','1','0'),
            ('0','0','1','0','1','0','1','0','1','0','1','1','0','0'),
            ('0','0','1','0','1','0','1','0','1','0','1','1','1','0'),
            ('0','0','1','0','1','0','1','0','1','1','0','0','0','0'),
            ('0','0','1','0','1','0','1','0','1','1','0','0','1','0'),
            ('0','0','1','0','1','0','1','0','1','1','0','1','0','0'),
            ('0','0','1','0','1','0','1','0','1','1','0','1','1','0'),
            ('0','0','1','0','1','0','1','0','1','1','1','0','0','0'),
            ('0','0','1','0','1','0','1','0','1','1','1','0','1','0'),
            ('0','0','1','0','1','0','1','0','1','1','1','1','0','0'),
            ('0','0','1','0','1','0','1','0','1','1','1','1','1','0'),
            ('0','0','1','0','1','0','1','1','0','0','0','0','0','0'),
            ('0','0','1','0','1','0','1','1','0','0','0','0','1','0'),
            ('0','0','1','0','1','0','1','1','0','0','0','1','0','0'),
            ('0','0','1','0','1','0','1','1','0','0','0','1','1','0'),
            ('0','0','1','0','1','0','1','1','0','0','1','0','0','0'),
            ('0','0','1','0','1','0','1','1','0','0','1','0','1','0'),
            ('0','0','1','0','1','0','1','1','0','0','1','1','0','0'),
            ('0','0','1','0','1','0','1','1','0','0','1','1','1','0'),
            ('0','0','1','0','1','0','1','1','0','1','0','0','0','0'),
            ('0','0','1','0','1','0','1','1','0','1','0','0','1','0'),
            ('0','0','1','0','1','0','1','1','0','1','0','1','0','0'),
            ('0','0','1','0','1','0','1','1','0','1','0','1','1','0'),
            ('0','0','1','0','1','0','1','1','0','1','1','0','0','0'),
            ('0','0','1','0','1','0','1','1','0','1','1','0','1','0'),
            ('0','0','1','0','1','0','1','1','0','1','1','1','0','0'),
            ('0','0','1','0','1','0','1','1','0','1','1','1','1','0'),
            ('0','0','1','0','1','0','1','1','1','0','0','0','0','0'),
            ('0','0','1','0','1','0','1','1','1','0','0','0','1','0'),
            ('0','0','1','0','1','0','1','1','1','0','0','1','0','0'),
            ('0','0','1','0','1','0','1','1','1','0','0','1','1','0'),
            ('0','0','1','0','1','0','1','1','1','0','1','0','0','0'),
            ('0','0','1','0','1','0','1','1','1','0','1','0','1','0'),
            ('0','0','1','0','1','0','1','1','1','0','1','1','0','0'),
            ('0','0','1','0','1','0','1','1','1','0','1','1','1','0'),
            ('0','0','1','0','1','0','1','1','1','1','0','0','0','0'),
            ('0','0','1','0','1','0','1','1','1','1','0','0','1','0'),
            ('0','0','1','0','1','0','1','1','1','1','0','1','0','0'),
            ('0','0','1','0','1','0','1','1','1','1','0','1','1','0'),
            ('0','0','1','0','1','0','1','1','1','1','1','0','0','0'),
            ('0','0','1','0','1','0','1','1','1','1','1','0','1','0'),
            ('0','0','1','0','1','0','1','1','1','1','1','1','0','0'),
            ('0','0','1','0','1','0','1','1','1','1','1','1','1','0'),
            ('0','0','1','0','1','1','0','0','0','0','0','0','0','0'),
            ('0','0','1','0','1','1','0','0','0','0','0','0','1','0'),
            ('0','0','1','0','1','1','0','0','0','0','0','1','0','0'),
            ('0','0','1','0','1','1','0','0','0','0','0','1','1','0'),
            ('0','0','1','0','1','1','0','0','0','0','1','0','0','0'),
            ('0','0','1','0','1','1','0','0','0','0','1','0','1','0'),
            ('0','0','1','0','1','1','0','0','0','0','1','1','0','0'),
            ('0','0','1','0','1','1','0','0','0','0','1','1','1','0'),
            ('0','0','1','0','1','1','0','0','0','1','0','0','0','0'),
            ('0','0','1','0','1','1','0','0','0','1','0','0','1','0'),
            ('0','0','1','0','1','1','0','0','0','1','0','1','0','0'),
            ('0','0','1','0','1','1','0','0','0','1','0','1','1','0'),
            ('0','0','1','0','1','1','0','0','0','1','1','0','0','0'),
            ('0','0','1','0','1','1','0','0','0','1','1','0','1','0'),
            ('0','0','1','0','1','1','0','0','0','1','1','1','0','0'),
            ('0','0','1','0','1','1','0','0','0','1','1','1','1','0'),
            ('0','0','1','0','1','1','0','0','1','0','0','0','0','0'),
            ('0','0','1','0','1','1','0','0','1','0','0','0','1','0'),
            ('0','0','1','0','1','1','0','0','1','0','0','1','0','0'),
            ('0','0','1','0','1','1','0','0','1','0','0','1','1','0'),
            ('0','0','1','0','1','1','0','0','1','0','1','0','0','0'),
            ('0','0','1','0','1','1','0','0','1','0','1','0','1','0'),
            ('0','0','1','0','1','1','0','0','1','0','1','1','0','0'),
            ('0','0','1','0','1','1','0','0','1','0','1','1','1','0'),
            ('0','0','1','0','1','1','0','0','1','1','0','0','0','0'),
            ('0','0','1','0','1','1','0','0','1','1','0','0','1','0'),
            ('0','0','1','0','1','1','0','0','1','1','0','1','0','0'),
            ('0','0','1','0','1','1','0','0','1','1','0','1','1','0'),
            ('0','0','1','0','1','1','0','0','1','1','1','0','0','0'),
            ('0','0','1','0','1','1','0','0','1','1','1','0','1','0'),
            ('0','0','1','0','1','1','0','0','1','1','1','1','0','0'),
            ('0','0','1','0','1','1','0','0','1','1','1','1','1','0'),
            ('0','0','1','0','1','1','0','1','0','0','0','0','0','0'),
            ('0','0','1','0','1','1','0','1','0','0','0','0','1','0'),
            ('0','0','1','0','1','1','0','1','0','0','0','1','0','0'),
            ('0','0','1','0','1','1','0','1','0','0','0','1','1','0'),
            ('0','0','1','0','1','1','0','1','0','0','1','0','0','0'),
            ('0','0','1','0','1','1','0','1','0','0','1','0','1','0'),
            ('0','0','1','0','1','1','0','1','0','0','1','1','0','0'),
            ('0','0','1','0','1','1','0','1','0','0','1','1','1','0'),
            ('0','0','1','0','1','1','0','1','0','1','0','0','0','0'),
            ('0','0','1','0','1','1','0','1','0','1','0','0','1','0'),
            ('0','0','1','0','1','1','0','1','0','1','0','1','0','0'),
            ('0','0','1','0','1','1','0','1','0','1','0','1','1','0'),
            ('0','0','1','0','1','1','0','1','0','1','1','0','0','0'),
            ('0','0','1','0','1','1','0','1','0','1','1','0','1','0'),
            ('0','0','1','0','1','1','0','1','0','1','1','1','0','0'),
            ('0','0','1','0','1','1','0','1','0','1','1','1','1','0'),
            ('0','0','1','0','1','1','0','1','1','0','0','0','0','0'),
            ('0','0','1','0','1','1','0','1','1','0','0','0','1','0'),
            ('0','0','1','0','1','1','0','1','1','0','0','1','0','0'),
            ('0','0','1','0','1','1','0','1','1','0','0','1','1','0'),
            ('0','0','1','0','1','1','0','1','1','0','1','0','0','0'),
            ('0','0','1','0','1','1','0','1','1','0','1','0','1','0'),
            ('0','0','1','0','1','1','0','1','1','0','1','1','0','0'),
            ('0','0','1','0','1','1','0','1','1','0','1','1','1','0'),
            ('0','0','1','0','1','1','0','1','1','1','0','0','0','0'),
            ('0','0','1','0','1','1','0','1','1','1','0','0','1','0'),
            ('0','0','1','0','1','1','0','1','1','1','0','1','0','0'),
            ('0','0','1','0','1','1','0','1','1','1','0','1','1','0'),
            ('0','0','1','0','1','1','0','1','1','1','1','0','0','0'),
            ('0','0','1','0','1','1','0','1','1','1','1','0','1','0'),
            ('0','0','1','0','1','1','0','1','1','1','1','1','0','0'),
            ('0','0','1','0','1','1','0','1','1','1','1','1','1','0'),
            ('0','0','1','0','1','1','1','0','0','0','0','0','0','0'),
            ('0','0','1','0','1','1','1','0','0','0','0','0','1','0'),
            ('0','0','1','0','1','1','1','0','0','0','0','1','0','0'),
            ('0','0','1','0','1','1','1','0','0','0','0','1','1','0'),
            ('0','0','1','0','1','1','1','0','0','0','1','0','0','0'),
            ('0','0','1','0','1','1','1','0','0','0','1','0','1','0'),
            ('0','0','1','0','1','1','1','0','0','0','1','1','0','0'),
            ('0','0','1','0','1','1','1','0','0','0','1','1','1','0'),
            ('0','0','1','0','1','1','1','0','0','1','0','0','0','0'),
            ('0','0','1','0','1','1','1','0','0','1','0','0','1','0'),
            ('0','0','1','0','1','1','1','0','0','1','0','1','0','0'),
            ('0','0','1','0','1','1','1','0','0','1','0','1','1','0'),
            ('0','0','1','0','1','1','1','0','0','1','1','0','0','0'),
            ('0','0','1','0','1','1','1','0','0','1','1','0','1','0'),
            ('0','0','1','0','1','1','1','0','0','1','1','1','0','0'),
            ('0','0','1','0','1','1','1','0','0','1','1','1','1','0'),
            ('0','0','1','0','1','1','1','0','1','0','0','0','0','0'),
            ('0','0','1','0','1','1','1','0','1','0','0','0','1','0'),
            ('0','0','1','0','1','1','1','0','1','0','0','1','0','0'),
            ('0','0','1','0','1','1','1','0','1','0','0','1','1','0'),
            ('0','0','1','0','1','1','1','0','1','0','1','0','0','0'),
            ('0','0','1','0','1','1','1','0','1','0','1','0','1','0'),
            ('0','0','1','0','1','1','1','0','1','0','1','1','0','0'),
            ('0','0','1','0','1','1','1','0','1','0','1','1','1','0'),
            ('0','0','1','0','1','1','1','0','1','1','0','0','0','0'),
            ('0','0','1','0','1','1','1','0','1','1','0','0','1','0'),
            ('0','0','1','0','1','1','1','0','1','1','0','1','0','0'),
            ('0','0','1','0','1','1','1','0','1','1','0','1','1','0'),
            ('0','0','1','0','1','1','1','0','1','1','1','0','0','0'),
            ('0','0','1','0','1','1','1','0','1','1','1','0','1','0'),
            ('0','0','1','0','1','1','1','0','1','1','1','1','0','0'),
            ('0','0','1','0','1','1','1','0','1','1','1','1','1','0'),
            ('0','0','1','0','1','1','1','1','0','0','0','0','0','0'),
            ('0','0','1','0','1','1','1','1','0','0','0','0','1','0'),
            ('0','0','1','0','1','1','1','1','0','0','0','1','0','0'),
            ('0','0','1','0','1','1','1','1','0','0','0','1','1','0'),
            ('0','0','1','0','1','1','1','1','0','0','1','0','0','0'),
            ('0','0','1','0','1','1','1','1','0','0','1','0','1','0'),
            ('0','0','1','0','1','1','1','1','0','0','1','1','0','0'),
            ('0','0','1','0','1','1','1','1','0','0','1','1','1','0'),
            ('0','0','1','0','1','1','1','1','0','1','0','0','0','0'),
            ('0','0','1','0','1','1','1','1','0','1','0','0','1','0'),
            ('0','0','1','0','1','1','1','1','0','1','0','1','0','0'),
            ('0','0','1','0','1','1','1','1','0','1','0','1','1','0'),
            ('0','0','1','0','1','1','1','1','0','1','1','0','0','0'),
            ('0','0','1','0','1','1','1','1','0','1','1','0','1','0'),
            ('0','0','1','0','1','1','1','1','0','1','1','1','0','0'),
            ('0','0','1','0','1','1','1','1','0','1','1','1','1','0'),
            ('0','0','1','0','1','1','1','1','1','0','0','0','0','0'),
            ('0','0','1','0','1','1','1','1','1','0','0','0','1','0'),
            ('0','0','1','0','1','1','1','1','1','0','0','1','0','0'),
            ('0','0','1','0','1','1','1','1','1','0','0','1','1','0'),
            ('0','0','1','0','1','1','1','1','1','0','1','0','0','0'),
            ('0','0','1','0','1','1','1','1','1','0','1','0','1','0'),
            ('0','0','1','0','1','1','1','1','1','0','1','1','0','0'),
            ('0','0','1','0','1','1','1','1','1','0','1','1','1','0'),
            ('0','0','1','0','1','1','1','1','1','1','0','0','0','0'),
            ('0','0','1','0','1','1','1','1','1','1','0','0','1','0'),
            ('0','0','1','0','1','1','1','1','1','1','0','1','0','0'),
            ('0','0','1','0','1','1','1','1','1','1','0','1','1','0'),
            ('0','0','1','0','1','1','1','1','1','1','1','0','0','0'),
            ('0','0','1','0','1','1','1','1','1','1','1','0','1','0'),
            ('0','0','1','0','1','1','1','1','1','1','1','1','0','0'),
            ('0','0','1','0','1','1','1','1','1','1','1','1','1','0'),
            ('0','0','1','1','0','0','0','0','0','0','0','0','0','0'),
            ('0','0','1','1','0','0','0','0','0','0','0','0','1','0'),
            ('0','0','1','1','0','0','0','0','0','0','0','1','0','0'),
            ('0','0','1','1','0','0','0','0','0','0','0','1','1','0'),
            ('0','0','1','1','0','0','0','0','0','0','1','0','0','0'),
            ('0','0','1','1','0','0','0','0','0','0','1','0','1','0'),
            ('0','0','1','1','0','0','0','0','0','0','1','1','0','0'),
            ('0','0','1','1','0','0','0','0','0','0','1','1','1','0'),
            ('0','0','1','1','0','0','0','0','0','1','0','0','0','0'),
            ('0','0','1','1','0','0','0','0','0','1','0','0','1','0'),
            ('0','0','1','1','0','0','0','0','0','1','0','1','0','0'),
            ('0','0','1','1','0','0','0','0','0','1','0','1','1','0'),
            ('0','0','1','1','0','0','0','0','0','1','1','0','0','0'),
            ('0','0','1','1','0','0','0','0','0','1','1','0','1','0'),
            ('0','0','1','1','0','0','0','0','0','1','1','1','0','0'),
            ('0','0','1','1','0','0','0','0','0','1','1','1','1','0'),
            ('0','0','1','1','0','0','0','0','1','0','0','0','0','0'),
            ('0','0','1','1','0','0','0','0','1','0','0','0','1','0'),
            ('0','0','1','1','0','0','0','0','1','0','0','1','0','0'),
            ('0','0','1','1','0','0','0','0','1','0','0','1','1','0'),
            ('0','0','1','1','0','0','0','0','1','0','1','0','0','0'),
            ('0','0','1','1','0','0','0','0','1','0','1','0','1','0'),
            ('0','0','1','1','0','0','0','0','1','0','1','1','0','0'),
            ('0','0','1','1','0','0','0','0','1','0','1','1','1','0'),
            ('0','0','1','1','0','0','0','0','1','1','0','0','0','0'),
            ('0','0','1','1','0','0','0','0','1','1','0','0','1','0'),
            ('0','0','1','1','0','0','0','0','1','1','0','1','0','0'),
            ('0','0','1','1','0','0','0','0','1','1','0','1','1','0'),
            ('0','0','1','1','0','0','0','0','1','1','1','0','0','0'),
            ('0','0','1','1','0','0','0','0','1','1','1','0','1','0'),
            ('0','0','1','1','0','0','0','0','1','1','1','1','0','0'),
            ('0','0','1','1','0','0','0','0','1','1','1','1','1','0'),
            ('0','0','1','1','0','0','0','1','0','0','0','0','0','0'),
            ('0','0','1','1','0','0','0','1','0','0','0','0','1','0'),
            ('0','0','1','1','0','0','0','1','0','0','0','1','0','0'),
            ('0','0','1','1','0','0','0','1','0','0','0','1','1','0'),
            ('0','0','1','1','0','0','0','1','0','0','1','0','0','0'),
            ('0','0','1','1','0','0','0','1','0','0','1','0','1','0'),
            ('0','0','1','1','0','0','0','1','0','0','1','1','0','0'),
            ('0','0','1','1','0','0','0','1','0','0','1','1','1','0'),
            ('0','0','1','1','0','0','0','1','0','1','0','0','0','0'),
            ('0','0','1','1','0','0','0','1','0','1','0','0','1','0'),
            ('0','0','1','1','0','0','0','1','0','1','0','1','0','0'),
            ('0','0','1','1','0','0','0','1','0','1','0','1','1','0'),
            ('0','0','1','1','0','0','0','1','0','1','1','0','0','0'),
            ('0','0','1','1','0','0','0','1','0','1','1','0','1','0'),
            ('0','0','1','1','0','0','0','1','0','1','1','1','0','0'),
            ('0','0','1','1','0','0','0','1','0','1','1','1','1','0'),
            ('0','0','1','1','0','0','0','1','1','0','0','0','0','0'),
            ('0','0','1','1','0','0','0','1','1','0','0','0','1','0'),
            ('0','0','1','1','0','0','0','1','1','0','0','1','0','0'),
            ('0','0','1','1','0','0','0','1','1','0','0','1','1','0'),
            ('0','0','1','1','0','0','0','1','1','0','1','0','0','0'),
            ('0','0','1','1','0','0','0','1','1','0','1','0','1','0'),
            ('0','0','1','1','0','0','0','1','1','0','1','1','0','0'),
            ('0','0','1','1','0','0','0','1','1','0','1','1','1','0'),
            ('0','0','1','1','0','0','0','1','1','1','0','0','0','0'),
            ('0','0','1','1','0','0','0','1','1','1','0','0','1','0'),
            ('0','0','1','1','0','0','0','1','1','1','0','1','0','0'),
            ('0','0','1','1','0','0','0','1','1','1','0','1','1','0'),
            ('0','0','1','1','0','0','0','1','1','1','1','0','0','0'),
            ('0','0','1','1','0','0','0','1','1','1','1','0','1','0'),
            ('0','0','1','1','0','0','0','1','1','1','1','1','0','0'),
            ('0','0','1','1','0','0','0','1','1','1','1','1','1','0'),
            ('0','0','1','1','0','0','1','0','0','0','0','0','0','0'),
            ('0','0','1','1','0','0','1','0','0','0','0','0','1','0'),
            ('0','0','1','1','0','0','1','0','0','0','0','1','0','0'),
            ('0','0','1','1','0','0','1','0','0','0','0','1','1','0'),
            ('0','0','1','1','0','0','1','0','0','0','1','0','0','0'),
            ('0','0','1','1','0','0','1','0','0','0','1','0','1','0'),
            ('0','0','1','1','0','0','1','0','0','0','1','1','0','0'),
            ('0','0','1','1','0','0','1','0','0','0','1','1','1','0'),
            ('0','0','1','1','0','0','1','0','0','1','0','0','0','0'),
            ('0','0','1','1','0','0','1','0','0','1','0','0','1','0'),
            ('0','0','1','1','0','0','1','0','0','1','0','1','0','0'),
            ('0','0','1','1','0','0','1','0','0','1','0','1','1','0'),
            ('0','0','1','1','0','0','1','0','0','1','1','0','0','0'),
            ('0','0','1','1','0','0','1','0','0','1','1','0','1','0'),
            ('0','0','1','1','0','0','1','0','0','1','1','1','0','0'),
            ('0','0','1','1','0','0','1','0','0','1','1','1','1','0'),
            ('0','0','1','1','0','0','1','0','1','0','0','0','0','0'),
            ('0','0','1','1','0','0','1','0','1','0','0','0','1','0'),
            ('0','0','1','1','0','0','1','0','1','0','0','1','0','0'),
            ('0','0','1','1','0','0','1','0','1','0','0','1','1','0'),
            ('0','0','1','1','0','0','1','0','1','0','1','0','0','0'),
            ('0','0','1','1','0','0','1','0','1','0','1','0','1','0'),
            ('0','0','1','1','0','0','1','0','1','0','1','1','0','0'),
            ('0','0','1','1','0','0','1','0','1','0','1','1','1','0'),
            ('0','0','1','1','0','0','1','0','1','1','0','0','0','0'),
            ('0','0','1','1','0','0','1','0','1','1','0','0','1','0'),
            ('0','0','1','1','0','0','1','0','1','1','0','1','0','0'),
            ('0','0','1','1','0','0','1','0','1','1','0','1','1','0'),
            ('0','0','1','1','0','0','1','0','1','1','1','0','0','0'),
            ('0','0','1','1','0','0','1','0','1','1','1','0','1','0'),
            ('0','0','1','1','0','0','1','0','1','1','1','1','0','0'),
            ('0','0','1','1','0','0','1','0','1','1','1','1','1','0'),
            ('0','0','1','1','0','0','1','1','0','0','0','0','0','0'),
            ('0','0','1','1','0','0','1','1','0','0','0','0','1','0'),
            ('0','0','1','1','0','0','1','1','0','0','0','1','0','0'),
            ('0','0','1','1','0','0','1','1','0','0','0','1','1','0'),
            ('0','0','1','1','0','0','1','1','0','0','1','0','0','0'),
            ('0','0','1','1','0','0','1','1','0','0','1','0','1','0'),
            ('0','0','1','1','0','0','1','1','0','0','1','1','0','0'),
            ('0','0','1','1','0','0','1','1','0','0','1','1','1','0'),
            ('0','0','1','1','0','0','1','1','0','1','0','0','0','0'),
            ('0','0','1','1','0','0','1','1','0','1','0','0','1','0'),
            ('0','0','1','1','0','0','1','1','0','1','0','1','0','0'),
            ('0','0','1','1','0','0','1','1','0','1','0','1','1','0'),
            ('0','0','1','1','0','0','1','1','0','1','1','0','0','0'),
            ('0','0','1','1','0','0','1','1','0','1','1','0','1','0'),
            ('0','0','1','1','0','0','1','1','0','1','1','1','0','0'),
            ('0','0','1','1','0','0','1','1','0','1','1','1','1','0'),
            ('0','0','1','1','0','0','1','1','1','0','0','0','0','0'),
            ('0','0','1','1','0','0','1','1','1','0','0','0','1','0'),
            ('0','0','1','1','0','0','1','1','1','0','0','1','0','0'),
            ('0','0','1','1','0','0','1','1','1','0','0','1','1','0'),
            ('0','0','1','1','0','0','1','1','1','0','1','0','0','0'),
            ('0','0','1','1','0','0','1','1','1','0','1','0','1','0'),
            ('0','0','1','1','0','0','1','1','1','0','1','1','0','0'),
            ('0','0','1','1','0','0','1','1','1','0','1','1','1','0'),
            ('0','0','1','1','0','0','1','1','1','1','0','0','0','0'),
            ('0','0','1','1','0','0','1','1','1','1','0','0','1','0'),
            ('0','0','1','1','0','0','1','1','1','1','0','1','0','0'),
            ('0','0','1','1','0','0','1','1','1','1','0','1','1','0'),
            ('0','0','1','1','0','0','1','1','1','1','1','0','0','0'),
            ('0','0','1','1','0','0','1','1','1','1','1','0','1','0'),
            ('0','0','1','1','0','0','1','1','1','1','1','1','0','0'),
            ('0','0','1','1','0','0','1','1','1','1','1','1','1','0'),
            ('0','0','1','1','0','1','0','0','0','0','0','0','0','0'),
            ('0','0','1','1','0','1','0','0','0','0','0','0','1','0'),
            ('0','0','1','1','0','1','0','0','0','0','0','1','0','0'),
            ('0','0','1','1','0','1','0','0','0','0','0','1','1','0'),
            ('0','0','1','1','0','1','0','0','0','0','1','0','0','0'),
            ('0','0','1','1','0','1','0','0','0','0','1','0','1','0'),
            ('0','0','1','1','0','1','0','0','0','0','1','1','0','0'),
            ('0','0','1','1','0','1','0','0','0','0','1','1','1','0'),
            ('0','0','1','1','0','1','0','0','0','1','0','0','0','0'),
            ('0','0','1','1','0','1','0','0','0','1','0','0','1','0'),
            ('0','0','1','1','0','1','0','0','0','1','0','1','0','0'),
            ('0','0','1','1','0','1','0','0','0','1','0','1','1','0'),
            ('0','0','1','1','0','1','0','0','0','1','1','0','0','0'),
            ('0','0','1','1','0','1','0','0','0','1','1','0','1','0'),
            ('0','0','1','1','0','1','0','0','0','1','1','1','0','0'),
            ('0','0','1','1','0','1','0','0','0','1','1','1','1','0'),
            ('0','0','1','1','0','1','0','0','1','0','0','0','0','0'),
            ('0','0','1','1','0','1','0','0','1','0','0','0','1','0'),
            ('0','0','1','1','0','1','0','0','1','0','0','1','0','0'),
            ('0','0','1','1','0','1','0','0','1','0','0','1','1','0'),
            ('0','0','1','1','0','1','0','0','1','0','1','0','0','0'),
            ('0','0','1','1','0','1','0','0','1','0','1','0','1','0'),
            ('0','0','1','1','0','1','0','0','1','0','1','1','0','0'),
            ('0','0','1','1','0','1','0','0','1','0','1','1','1','0'),
            ('0','0','1','1','0','1','0','0','1','1','0','0','0','0'),
            ('0','0','1','1','0','1','0','0','1','1','0','0','1','0'),
            ('0','0','1','1','0','1','0','0','1','1','0','1','0','0'),
            ('0','0','1','1','0','1','0','0','1','1','0','1','1','0'),
            ('0','0','1','1','0','1','0','0','1','1','1','0','0','0'),
            ('0','0','1','1','0','1','0','0','1','1','1','0','1','0'),
            ('0','0','1','1','0','1','0','0','1','1','1','1','0','0'),
            ('0','0','1','1','0','1','0','0','1','1','1','1','1','0'),
            ('0','0','1','1','0','1','0','1','0','0','0','0','0','0'),
            ('0','0','1','1','0','1','0','1','0','0','0','0','1','0'),
            ('0','0','1','1','0','1','0','1','0','0','0','1','0','0'),
            ('0','0','1','1','0','1','0','1','0','0','0','1','1','0'),
            ('0','0','1','1','0','1','0','1','0','0','1','0','0','0'),
            ('0','0','1','1','0','1','0','1','0','0','1','0','1','0'),
            ('0','0','1','1','0','1','0','1','0','0','1','1','0','0'),
            ('0','0','1','1','0','1','0','1','0','0','1','1','1','0'),
            ('0','0','1','1','0','1','0','1','0','1','0','0','0','0'),
            ('0','0','1','1','0','1','0','1','0','1','0','0','1','0'),
            ('0','0','1','1','0','1','0','1','0','1','0','1','0','0'),
            ('0','0','1','1','0','1','0','1','0','1','0','1','1','0'),
            ('0','0','1','1','0','1','0','1','0','1','1','0','0','0'),
            ('0','0','1','1','0','1','0','1','0','1','1','0','1','0'),
            ('0','0','1','1','0','1','0','1','0','1','1','1','0','0'),
            ('0','0','1','1','0','1','0','1','0','1','1','1','1','0'),
            ('0','0','1','1','0','1','0','1','1','0','0','0','0','0'),
            ('0','0','1','1','0','1','0','1','1','0','0','0','1','0'),
            ('0','0','1','1','0','1','0','1','1','0','0','1','0','0'),
            ('0','0','1','1','0','1','0','1','1','0','0','1','1','0'),
            ('0','0','1','1','0','1','0','1','1','0','1','0','0','0'),
            ('0','0','1','1','0','1','0','1','1','0','1','0','1','0'),
            ('0','0','1','1','0','1','0','1','1','0','1','1','0','0'),
            ('0','0','1','1','0','1','0','1','1','0','1','1','1','0'),
            ('0','0','1','1','0','1','0','1','1','1','0','0','0','0'),
            ('0','0','1','1','0','1','0','1','1','1','0','0','1','0'),
            ('0','0','1','1','0','1','0','1','1','1','0','1','0','0'),
            ('0','0','1','1','0','1','0','1','1','1','0','1','1','0'),
            ('0','0','1','1','0','1','0','1','1','1','1','0','0','0'),
            ('0','0','1','1','0','1','0','1','1','1','1','0','1','0'),
            ('0','0','1','1','0','1','0','1','1','1','1','1','0','0'),
            ('0','0','1','1','0','1','0','1','1','1','1','1','1','0'),
            ('0','0','1','1','0','1','1','0','0','0','0','0','0','0'),
            ('0','0','1','1','0','1','1','0','0','0','0','0','1','0'),
            ('0','0','1','1','0','1','1','0','0','0','0','1','0','0'),
            ('0','0','1','1','0','1','1','0','0','0','0','1','1','0'),
            ('0','0','1','1','0','1','1','0','0','0','1','0','0','0'),
            ('0','0','1','1','0','1','1','0','0','0','1','0','1','0'),
            ('0','0','1','1','0','1','1','0','0','0','1','1','0','0'),
            ('0','0','1','1','0','1','1','0','0','0','1','1','1','0'),
            ('0','0','1','1','0','1','1','0','0','1','0','0','0','0'),
            ('0','0','1','1','0','1','1','0','0','1','0','0','1','0'),
            ('0','0','1','1','0','1','1','0','0','1','0','1','0','0'),
            ('0','0','1','1','0','1','1','0','0','1','0','1','1','0'),
            ('0','0','1','1','0','1','1','0','0','1','1','0','0','0'),
            ('0','0','1','1','0','1','1','0','0','1','1','0','1','0'),
            ('0','0','1','1','0','1','1','0','0','1','1','1','0','0'),
            ('0','0','1','1','0','1','1','0','0','1','1','1','1','0'),
            ('0','0','1','1','0','1','1','0','1','0','0','0','0','0'),
            ('0','0','1','1','0','1','1','0','1','0','0','0','1','0'),
            ('0','0','1','1','0','1','1','0','1','0','0','1','0','0'),
            ('0','0','1','1','0','1','1','0','1','0','0','1','1','0'),
            ('0','0','1','1','0','1','1','0','1','0','1','0','0','0'),
            ('0','0','1','1','0','1','1','0','1','0','1','0','1','0'),
            ('0','0','1','1','0','1','1','0','1','0','1','1','0','0'),
            ('0','0','1','1','0','1','1','0','1','0','1','1','1','0'),
            ('0','0','1','1','0','1','1','0','1','1','0','0','0','0'),
            ('0','0','1','1','0','1','1','0','1','1','0','0','1','0'),
            ('0','0','1','1','0','1','1','0','1','1','0','1','0','0'),
            ('0','0','1','1','0','1','1','0','1','1','0','1','1','0'),
            ('0','0','1','1','0','1','1','0','1','1','1','0','0','0'),
            ('0','0','1','1','0','1','1','0','1','1','1','0','1','0'),
            ('0','0','1','1','0','1','1','0','1','1','1','1','0','0'),
            ('0','0','1','1','0','1','1','0','1','1','1','1','1','0'),
            ('0','0','1','1','0','1','1','1','0','0','0','0','0','0'),
            ('0','0','1','1','0','1','1','1','0','0','0','0','1','0'),
            ('0','0','1','1','0','1','1','1','0','0','0','1','0','0'),
            ('0','0','1','1','0','1','1','1','0','0','0','1','1','0'),
            ('0','0','1','1','0','1','1','1','0','0','1','0','0','0'),
            ('0','0','1','1','0','1','1','1','0','0','1','0','1','0'),
            ('0','0','1','1','0','1','1','1','0','0','1','1','0','0'),
            ('0','0','1','1','0','1','1','1','0','0','1','1','1','0'),
            ('0','0','1','1','0','1','1','1','0','1','0','0','0','0'),
            ('0','0','1','1','0','1','1','1','0','1','0','0','1','0'),
            ('0','0','1','1','0','1','1','1','0','1','0','1','0','0'),
            ('0','0','1','1','0','1','1','1','0','1','0','1','1','0'),
            ('0','0','1','1','0','1','1','1','0','1','1','0','0','0'),
            ('0','0','1','1','0','1','1','1','0','1','1','0','1','0'),
            ('0','0','1','1','0','1','1','1','0','1','1','1','0','0'),
            ('0','0','1','1','0','1','1','1','0','1','1','1','1','0'),
            ('0','0','1','1','0','1','1','1','1','0','0','0','0','0'),
            ('0','0','1','1','0','1','1','1','1','0','0','0','1','0'),
            ('0','0','1','1','0','1','1','1','1','0','0','1','0','0'),
            ('0','0','1','1','0','1','1','1','1','0','0','1','1','0'),
            ('0','0','1','1','0','1','1','1','1','0','1','0','0','0'),
            ('0','0','1','1','0','1','1','1','1','0','1','0','1','0'),
            ('0','0','1','1','0','1','1','1','1','0','1','1','0','0'),
            ('0','0','1','1','0','1','1','1','1','0','1','1','1','0'),
            ('0','0','1','1','0','1','1','1','1','1','0','0','0','0'),
            ('0','0','1','1','0','1','1','1','1','1','0','0','1','0'),
            ('0','0','1','1','0','1','1','1','1','1','0','1','0','0'),
            ('0','0','1','1','0','1','1','1','1','1','0','1','1','0'),
            ('0','0','1','1','0','1','1','1','1','1','1','0','0','0'),
            ('0','0','1','1','0','1','1','1','1','1','1','0','1','0'),
            ('0','0','1','1','0','1','1','1','1','1','1','1','0','0'),
            ('0','0','1','1','0','1','1','1','1','1','1','1','1','0'),
            ('0','0','1','1','1','0','0','0','0','0','0','0','0','0'),
            ('0','0','1','1','1','0','0','0','0','0','0','0','1','0'),
            ('0','0','1','1','1','0','0','0','0','0','0','1','0','0'),
            ('0','0','1','1','1','0','0','0','0','0','0','1','1','0'),
            ('0','0','1','1','1','0','0','0','0','0','1','0','0','0'),
            ('0','0','1','1','1','0','0','0','0','0','1','0','1','0'),
            ('0','0','1','1','1','0','0','0','0','0','1','1','0','0'),
            ('0','0','1','1','1','0','0','0','0','0','1','1','1','0'),
            ('0','0','1','1','1','0','0','0','0','1','0','0','0','0'),
            ('0','0','1','1','1','0','0','0','0','1','0','0','1','0'),
            ('0','0','1','1','1','0','0','0','0','1','0','1','0','0'),
            ('0','0','1','1','1','0','0','0','0','1','0','1','1','0'),
            ('0','0','1','1','1','0','0','0','0','1','1','0','0','0'),
            ('0','0','1','1','1','0','0','0','0','1','1','0','1','0'),
            ('0','0','1','1','1','0','0','0','0','1','1','1','0','0'),
            ('0','0','1','1','1','0','0','0','0','1','1','1','1','0'),
            ('0','0','1','1','1','0','0','0','1','0','0','0','0','0'),
            ('0','0','1','1','1','0','0','0','1','0','0','0','1','0'),
            ('0','0','1','1','1','0','0','0','1','0','0','1','0','0'),
            ('0','0','1','1','1','0','0','0','1','0','0','1','1','0'),
            ('0','0','1','1','1','0','0','0','1','0','1','0','0','0'),
            ('0','0','1','1','1','0','0','0','1','0','1','0','1','0'),
            ('0','0','1','1','1','0','0','0','1','0','1','1','0','0'),
            ('0','0','1','1','1','0','0','0','1','0','1','1','1','0'),
            ('0','0','1','1','1','0','0','0','1','1','0','0','0','0'),
            ('0','0','1','1','1','0','0','0','1','1','0','0','1','0'),
            ('0','0','1','1','1','0','0','0','1','1','0','1','0','0'),
            ('0','0','1','1','1','0','0','0','1','1','0','1','1','0'),
            ('0','0','1','1','1','0','0','0','1','1','1','0','0','0'),
            ('0','0','1','1','1','0','0','0','1','1','1','0','1','0'),
            ('0','0','1','1','1','0','0','0','1','1','1','1','0','0'),
            ('0','0','1','1','1','0','0','0','1','1','1','1','1','0'),
            ('0','0','1','1','1','0','0','1','0','0','0','0','0','0'),
            ('0','0','1','1','1','0','0','1','0','0','0','0','1','0'),
            ('0','0','1','1','1','0','0','1','0','0','0','1','0','0'),
            ('0','0','1','1','1','0','0','1','0','0','0','1','1','0'),
            ('0','0','1','1','1','0','0','1','0','0','1','0','0','0'),
            ('0','0','1','1','1','0','0','1','0','0','1','0','1','0'),
            ('0','0','1','1','1','0','0','1','0','0','1','1','0','0'),
            ('0','0','1','1','1','0','0','1','0','0','1','1','1','0'),
            ('0','0','1','1','1','0','0','1','0','1','0','0','0','0'),
            ('0','0','1','1','1','0','0','1','0','1','0','0','1','0'),
            ('0','0','1','1','1','0','0','1','0','1','0','1','0','0'),
            ('0','0','1','1','1','0','0','1','0','1','0','1','1','0'),
            ('0','0','1','1','1','0','0','1','0','1','1','0','0','0'),
            ('0','0','1','1','1','0','0','1','0','1','1','0','1','0'),
            ('0','0','1','1','1','0','0','1','0','1','1','1','0','0'),
            ('0','0','1','1','1','0','0','1','0','1','1','1','1','0'),
            ('0','0','1','1','1','0','0','1','1','0','0','0','0','0'),
            ('0','0','1','1','1','0','0','1','1','0','0','0','1','0'),
            ('0','0','1','1','1','0','0','1','1','0','0','1','0','0'),
            ('0','0','1','1','1','0','0','1','1','0','0','1','1','0'),
            ('0','0','1','1','1','0','0','1','1','0','1','0','0','0'),
            ('0','0','1','1','1','0','0','1','1','0','1','0','1','0'),
            ('0','0','1','1','1','0','0','1','1','0','1','1','0','0'),
            ('0','0','1','1','1','0','0','1','1','0','1','1','1','0'),
            ('0','0','1','1','1','0','0','1','1','1','0','0','0','0'),
            ('0','0','1','1','1','0','0','1','1','1','0','0','1','0'),
            ('0','0','1','1','1','0','0','1','1','1','0','1','0','0'),
            ('0','0','1','1','1','0','0','1','1','1','0','1','1','0'),
            ('0','0','1','1','1','0','0','1','1','1','1','0','0','0'),
            ('0','0','1','1','1','0','0','1','1','1','1','0','1','0'),
            ('0','0','1','1','1','0','0','1','1','1','1','1','0','0'),
            ('0','0','1','1','1','0','0','1','1','1','1','1','1','0'),
            ('0','0','1','1','1','0','1','0','0','0','0','0','0','0'),
            ('0','0','1','1','1','0','1','0','0','0','0','0','1','0'),
            ('0','0','1','1','1','0','1','0','0','0','0','1','0','0'),
            ('0','0','1','1','1','0','1','0','0','0','0','1','1','0'),
            ('0','0','1','1','1','0','1','0','0','0','1','0','0','0'),
            ('0','0','1','1','1','0','1','0','0','0','1','0','1','0'),
            ('0','0','1','1','1','0','1','0','0','0','1','1','0','0'),
            ('0','0','1','1','1','0','1','0','0','0','1','1','1','0'),
            ('0','0','1','1','1','0','1','0','0','1','0','0','0','0'),
            ('0','0','1','1','1','0','1','0','0','1','0','0','1','0'),
            ('0','0','1','1','1','0','1','0','0','1','0','1','0','0'),
            ('0','0','1','1','1','0','1','0','0','1','0','1','1','0'),
            ('0','0','1','1','1','0','1','0','0','1','1','0','0','0'),
            ('0','0','1','1','1','0','1','0','0','1','1','0','1','0'),
            ('0','0','1','1','1','0','1','0','0','1','1','1','0','0'),
            ('0','0','1','1','1','0','1','0','0','1','1','1','1','0'),
            ('0','0','1','1','1','0','1','0','1','0','0','0','0','0'),
            ('0','0','1','1','1','0','1','0','1','0','0','0','1','0'),
            ('0','0','1','1','1','0','1','0','1','0','0','1','0','0'),
            ('0','0','1','1','1','0','1','0','1','0','0','1','1','0'),
            ('0','0','1','1','1','0','1','0','1','0','1','0','0','0'),
            ('0','0','1','1','1','0','1','0','1','0','1','0','1','0'),
            ('0','0','1','1','1','0','1','0','1','0','1','1','0','0'),
            ('0','0','1','1','1','0','1','0','1','0','1','1','1','0'),
            ('0','0','1','1','1','0','1','0','1','1','0','0','0','0'),
            ('0','0','1','1','1','0','1','0','1','1','0','0','1','0'),
            ('0','0','1','1','1','0','1','0','1','1','0','1','0','0'),
            ('0','0','1','1','1','0','1','0','1','1','0','1','1','0'),
            ('0','0','1','1','1','0','1','0','1','1','1','0','0','0'),
            ('0','0','1','1','1','0','1','0','1','1','1','0','1','0'),
            ('0','0','1','1','1','0','1','0','1','1','1','1','0','0'),
            ('0','0','1','1','1','0','1','0','1','1','1','1','1','0'),
            ('0','0','1','1','1','0','1','1','0','0','0','0','0','0'),
            ('0','0','1','1','1','0','1','1','0','0','0','0','1','0'),
            ('0','0','1','1','1','0','1','1','0','0','0','1','0','0'),
            ('0','0','1','1','1','0','1','1','0','0','0','1','1','0'),
            ('0','0','1','1','1','0','1','1','0','0','1','0','0','0'),
            ('0','0','1','1','1','0','1','1','0','0','1','0','1','0'),
            ('0','0','1','1','1','0','1','1','0','0','1','1','0','0'),
            ('0','0','1','1','1','0','1','1','0','0','1','1','1','0'),
            ('0','0','1','1','1','0','1','1','0','1','0','0','0','0'),
            ('0','0','1','1','1','0','1','1','0','1','0','0','1','0'),
            ('0','0','1','1','1','0','1','1','0','1','0','1','0','0'),
            ('0','0','1','1','1','0','1','1','0','1','0','1','1','0'),
            ('0','0','1','1','1','0','1','1','0','1','1','0','0','0'),
            ('0','0','1','1','1','0','1','1','0','1','1','0','1','0'),
            ('0','0','1','1','1','0','1','1','0','1','1','1','0','0'),
            ('0','0','1','1','1','0','1','1','0','1','1','1','1','0'),
            ('0','0','1','1','1','0','1','1','1','0','0','0','0','0'),
            ('0','0','1','1','1','0','1','1','1','0','0','0','1','0'),
            ('0','0','1','1','1','0','1','1','1','0','0','1','0','0'),
            ('0','0','1','1','1','0','1','1','1','0','0','1','1','0'),
            ('0','0','1','1','1','0','1','1','1','0','1','0','0','0'),
            ('0','0','1','1','1','0','1','1','1','0','1','0','1','0'),
            ('0','0','1','1','1','0','1','1','1','0','1','1','0','0'),
            ('0','0','1','1','1','0','1','1','1','0','1','1','1','0'),
            ('0','0','1','1','1','0','1','1','1','1','0','0','0','0'),
            ('0','0','1','1','1','0','1','1','1','1','0','0','1','0'),
            ('0','0','1','1','1','0','1','1','1','1','0','1','0','0'),
            ('0','0','1','1','1','0','1','1','1','1','0','1','1','0'),
            ('0','0','1','1','1','0','1','1','1','1','1','0','0','0'),
            ('0','0','1','1','1','0','1','1','1','1','1','0','1','0'),
            ('0','0','1','1','1','0','1','1','1','1','1','1','0','0'),
            ('0','0','1','1','1','0','1','1','1','1','1','1','1','0'),
            ('0','0','1','1','1','1','0','0','0','0','0','0','0','0'),
            ('0','0','1','1','1','1','0','0','0','0','0','0','1','0'),
            ('0','0','1','1','1','1','0','0','0','0','0','1','0','0'),
            ('0','0','1','1','1','1','0','0','0','0','0','1','1','0'),
            ('0','0','1','1','1','1','0','0','0','0','1','0','0','0'),
            ('0','0','1','1','1','1','0','0','0','0','1','0','1','0'),
            ('0','0','1','1','1','1','0','0','0','0','1','1','0','0'),
            ('0','0','1','1','1','1','0','0','0','0','1','1','1','0'),
            ('0','0','1','1','1','1','0','0','0','1','0','0','0','0'),
            ('0','0','1','1','1','1','0','0','0','1','0','0','1','0'),
            ('0','0','1','1','1','1','0','0','0','1','0','1','0','0'),
            ('0','0','1','1','1','1','0','0','0','1','0','1','1','0'),
            ('0','0','1','1','1','1','0','0','0','1','1','0','0','0'),
            ('0','0','1','1','1','1','0','0','0','1','1','0','1','0'),
            ('0','0','1','1','1','1','0','0','0','1','1','1','0','0'),
            ('0','0','1','1','1','1','0','0','0','1','1','1','1','0'),
            ('0','0','1','1','1','1','0','0','1','0','0','0','0','0'),
            ('0','0','1','1','1','1','0','0','1','0','0','0','1','0'),
            ('0','0','1','1','1','1','0','0','1','0','0','1','0','0'),
            ('0','0','1','1','1','1','0','0','1','0','0','1','1','0'),
            ('0','0','1','1','1','1','0','0','1','0','1','0','0','0'),
            ('0','0','1','1','1','1','0','0','1','0','1','0','1','0'),
            ('0','0','1','1','1','1','0','0','1','0','1','1','0','0'),
            ('0','0','1','1','1','1','0','0','1','0','1','1','1','0'),
            ('0','0','1','1','1','1','0','0','1','1','0','0','0','0'),
            ('0','0','1','1','1','1','0','0','1','1','0','0','1','0'),
            ('0','0','1','1','1','1','0','0','1','1','0','1','0','0'),
            ('0','0','1','1','1','1','0','0','1','1','0','1','1','0'),
            ('0','0','1','1','1','1','0','0','1','1','1','0','0','0'),
            ('0','0','1','1','1','1','0','0','1','1','1','0','1','0'),
            ('0','0','1','1','1','1','0','0','1','1','1','1','0','0'),
            ('0','0','1','1','1','1','0','0','1','1','1','1','1','0'),
            ('0','0','1','1','1','1','0','1','0','0','0','0','0','0'),
            ('0','0','1','1','1','1','0','1','0','0','0','0','1','0'),
            ('0','0','1','1','1','1','0','1','0','0','0','1','0','0'),
            ('0','0','1','1','1','1','0','1','0','0','0','1','1','0'),
            ('0','0','1','1','1','1','0','1','0','0','1','0','0','0'),
            ('0','0','1','1','1','1','0','1','0','0','1','0','1','0'),
            ('0','0','1','1','1','1','0','1','0','0','1','1','0','0'),
            ('0','0','1','1','1','1','0','1','0','0','1','1','1','0'),
            ('0','0','1','1','1','1','0','1','0','1','0','0','0','0'),
            ('0','0','1','1','1','1','0','1','0','1','0','0','1','0'),
            ('0','0','1','1','1','1','0','1','0','1','0','1','0','0'),
            ('0','0','1','1','1','1','0','1','0','1','0','1','1','0'),
            ('0','0','1','1','1','1','0','1','0','1','1','0','0','0'),
            ('0','0','1','1','1','1','0','1','0','1','1','0','1','0'),
            ('0','0','1','1','1','1','0','1','0','1','1','1','0','0'),
            ('0','0','1','1','1','1','0','1','0','1','1','1','1','0'),
            ('0','0','1','1','1','1','0','1','1','0','0','0','0','0'),
            ('0','0','1','1','1','1','0','1','1','0','0','0','1','0'),
            ('0','0','1','1','1','1','0','1','1','0','0','1','0','0'),
            ('0','0','1','1','1','1','0','1','1','0','0','1','1','0'),
            ('0','0','1','1','1','1','0','1','1','0','1','0','0','0'),
            ('0','0','1','1','1','1','0','1','1','0','1','0','1','0'),
            ('0','0','1','1','1','1','0','1','1','0','1','1','0','0'),
            ('0','0','1','1','1','1','0','1','1','0','1','1','1','0'),
            ('0','0','1','1','1','1','0','1','1','1','0','0','0','0'),
            ('0','0','1','1','1','1','0','1','1','1','0','0','1','0'),
            ('0','0','1','1','1','1','0','1','1','1','0','1','0','0'),
            ('0','0','1','1','1','1','0','1','1','1','0','1','1','0'),
            ('0','0','1','1','1','1','0','1','1','1','1','0','0','0'),
            ('0','0','1','1','1','1','0','1','1','1','1','0','1','0'),
            ('0','0','1','1','1','1','0','1','1','1','1','1','0','0'),
            ('0','0','1','1','1','1','0','1','1','1','1','1','1','0'),
            ('0','0','1','1','1','1','1','0','0','0','0','0','0','0'),
            ('0','0','1','1','1','1','1','0','0','0','0','0','1','0'),
            ('0','0','1','1','1','1','1','0','0','0','0','1','0','0'),
            ('0','0','1','1','1','1','1','0','0','0','0','1','1','0'),
            ('0','0','1','1','1','1','1','0','0','0','1','0','0','0'),
            ('0','0','1','1','1','1','1','0','0','0','1','0','1','0'),
            ('0','0','1','1','1','1','1','0','0','0','1','1','0','0'),
            ('0','0','1','1','1','1','1','0','0','0','1','1','1','0'),
            ('0','0','1','1','1','1','1','0','0','1','0','0','0','0'),
            ('0','0','1','1','1','1','1','0','0','1','0','0','1','0'),
            ('0','0','1','1','1','1','1','0','0','1','0','1','0','0'),
            ('0','0','1','1','1','1','1','0','0','1','0','1','1','0'),
            ('0','0','1','1','1','1','1','0','0','1','1','0','0','0'),
            ('0','0','1','1','1','1','1','0','0','1','1','0','1','0'),
            ('0','0','1','1','1','1','1','0','0','1','1','1','0','0'),
            ('0','0','1','1','1','1','1','0','0','1','1','1','1','0'),
            ('0','0','1','1','1','1','1','0','1','0','0','0','0','0'),
            ('0','0','1','1','1','1','1','0','1','0','0','0','1','0'),
            ('0','0','1','1','1','1','1','0','1','0','0','1','0','0'),
            ('0','0','1','1','1','1','1','0','1','0','0','1','1','0'),
            ('0','0','1','1','1','1','1','0','1','0','1','0','0','0'),
            ('0','0','1','1','1','1','1','0','1','0','1','0','1','0'),
            ('0','0','1','1','1','1','1','0','1','0','1','1','0','0'),
            ('0','0','1','1','1','1','1','0','1','0','1','1','1','0'),
            ('0','0','1','1','1','1','1','0','1','1','0','0','0','0'),
            ('0','0','1','1','1','1','1','0','1','1','0','0','1','0'),
            ('0','0','1','1','1','1','1','0','1','1','0','1','0','0'),
            ('0','0','1','1','1','1','1','0','1','1','0','1','1','0'),
            ('0','0','1','1','1','1','1','0','1','1','1','0','0','0'),
            ('0','0','1','1','1','1','1','0','1','1','1','0','1','0'),
            ('0','0','1','1','1','1','1','0','1','1','1','1','0','0'),
            ('0','0','1','1','1','1','1','0','1','1','1','1','1','0'),
            ('0','0','1','1','1','1','1','1','0','0','0','0','0','0'),
            ('0','0','1','1','1','1','1','1','0','0','0','0','1','0'),
            ('0','0','1','1','1','1','1','1','0','0','0','1','0','0'),
            ('0','0','1','1','1','1','1','1','0','0','0','1','1','0'),
            ('0','0','1','1','1','1','1','1','0','0','1','0','0','0'),
            ('0','0','1','1','1','1','1','1','0','0','1','0','1','0'),
            ('0','0','1','1','1','1','1','1','0','0','1','1','0','0'),
            ('0','0','1','1','1','1','1','1','0','0','1','1','1','0'),
            ('0','0','1','1','1','1','1','1','0','1','0','0','0','0'),
            ('0','0','1','1','1','1','1','1','0','1','0','0','1','0'),
            ('0','0','1','1','1','1','1','1','0','1','0','1','0','0'),
            ('0','0','1','1','1','1','1','1','0','1','0','1','1','0'),
            ('0','0','1','1','1','1','1','1','0','1','1','0','0','0'),
            ('0','0','1','1','1','1','1','1','0','1','1','0','1','0'),
            ('0','0','1','1','1','1','1','1','0','1','1','1','0','0'),
            ('0','0','1','1','1','1','1','1','0','1','1','1','1','0'),
            ('0','0','1','1','1','1','1','1','1','0','0','0','0','0'),
            ('0','0','1','1','1','1','1','1','1','0','0','0','1','0'),
            ('0','0','1','1','1','1','1','1','1','0','0','1','0','0'),
            ('0','0','1','1','1','1','1','1','1','0','0','1','1','0'),
            ('0','0','1','1','1','1','1','1','1','0','1','0','0','0'),
            ('0','0','1','1','1','1','1','1','1','0','1','0','1','0'),
            ('0','0','1','1','1','1','1','1','1','0','1','1','0','0'),
            ('0','0','1','1','1','1','1','1','1','0','1','1','1','0'),
            ('0','0','1','1','1','1','1','1','1','1','0','0','0','0'),
            ('0','0','1','1','1','1','1','1','1','1','0','0','1','0'),
            ('0','0','1','1','1','1','1','1','1','1','0','1','0','0'),
            ('0','0','1','1','1','1','1','1','1','1','0','1','1','0'),
            ('0','0','1','1','1','1','1','1','1','1','1','0','0','0'),
            ('0','0','1','1','1','1','1','1','1','1','1','0','1','0'),
            ('0','0','1','1','1','1','1','1','1','1','1','1','0','0'),
            ('0','0','1','1','1','1','1','1','1','1','1','1','1','0'),
            ('0','1','0','0','0','0','0','0','0','0','0','0','0','0'),
            ('0','1','0','0','0','0','0','0','0','0','0','0','1','0'),
            ('0','1','0','0','0','0','0','0','0','0','0','1','0','0'),
            ('0','1','0','0','0','0','0','0','0','0','0','1','1','0'),
            ('0','1','0','0','0','0','0','0','0','0','1','0','0','0'),
            ('0','1','0','0','0','0','0','0','0','0','1','0','1','0'),
            ('0','1','0','0','0','0','0','0','0','0','1','1','0','0'),
            ('0','1','0','0','0','0','0','0','0','0','1','1','1','0'),
            ('0','1','0','0','0','0','0','0','0','1','0','0','0','0'),
            ('0','1','0','0','0','0','0','0','0','1','0','0','1','0'),
            ('0','1','0','0','0','0','0','0','0','1','0','1','0','0'),
            ('0','1','0','0','0','0','0','0','0','1','0','1','1','0'),
            ('0','1','0','0','0','0','0','0','0','1','1','0','0','0'),
            ('0','1','0','0','0','0','0','0','0','1','1','0','1','0'),
            ('0','1','0','0','0','0','0','0','0','1','1','1','0','0'),
            ('0','1','0','0','0','0','0','0','0','1','1','1','1','0'),
            ('0','1','0','0','0','0','0','0','1','0','0','0','0','0'),
            ('0','1','0','0','0','0','0','0','1','0','0','0','1','0'),
            ('0','1','0','0','0','0','0','0','1','0','0','1','0','0'),
            ('0','1','0','0','0','0','0','0','1','0','0','1','1','0'),
            ('0','1','0','0','0','0','0','0','1','0','1','0','0','0'),
            ('0','1','0','0','0','0','0','0','1','0','1','0','1','0'),
            ('0','1','0','0','0','0','0','0','1','0','1','1','0','0'),
            ('0','1','0','0','0','0','0','0','1','0','1','1','1','0'),
            ('0','1','0','0','0','0','0','0','1','1','0','0','0','0'),
            ('0','1','0','0','0','0','0','0','1','1','0','0','1','0'),
            ('0','1','0','0','0','0','0','0','1','1','0','1','0','0'),
            ('0','1','0','0','0','0','0','0','1','1','0','1','1','0'),
            ('0','1','0','0','0','0','0','0','1','1','1','0','0','0'),
            ('0','1','0','0','0','0','0','0','1','1','1','0','1','0'),
            ('0','1','0','0','0','0','0','0','1','1','1','1','0','0'),
            ('0','1','0','0','0','0','0','0','1','1','1','1','1','0'),
            ('0','1','0','0','0','0','0','1','0','0','0','0','0','0'),
            ('0','1','0','0','0','0','0','1','0','0','0','0','1','0'),
            ('0','1','0','0','0','0','0','1','0','0','0','1','0','0'),
            ('0','1','0','0','0','0','0','1','0','0','0','1','1','0'),
            ('0','1','0','0','0','0','0','1','0','0','1','0','0','0'),
            ('0','1','0','0','0','0','0','1','0','0','1','0','1','0'),
            ('0','1','0','0','0','0','0','1','0','0','1','1','0','0'),
            ('0','1','0','0','0','0','0','1','0','0','1','1','1','0'),
            ('0','1','0','0','0','0','0','1','0','1','0','0','0','0'),
            ('0','1','0','0','0','0','0','1','0','1','0','0','1','0'),
            ('0','1','0','0','0','0','0','1','0','1','0','1','0','0'),
            ('0','1','0','0','0','0','0','1','0','1','0','1','1','0'),
            ('0','1','0','0','0','0','0','1','0','1','1','0','0','0'),
            ('0','1','0','0','0','0','0','1','0','1','1','0','1','0'),
            ('0','1','0','0','0','0','0','1','0','1','1','1','0','0'),
            ('0','1','0','0','0','0','0','1','0','1','1','1','1','0'),
            ('0','1','0','0','0','0','0','1','1','0','0','0','0','0'),
            ('0','1','0','0','0','0','0','1','1','0','0','0','1','0'),
            ('0','1','0','0','0','0','0','1','1','0','0','1','0','0'),
            ('0','1','0','0','0','0','0','1','1','0','0','1','1','0'),
            ('0','1','0','0','0','0','0','1','1','0','1','0','0','0'),
            ('0','1','0','0','0','0','0','1','1','0','1','0','1','0'),
            ('0','1','0','0','0','0','0','1','1','0','1','1','0','0'),
            ('0','1','0','0','0','0','0','1','1','0','1','1','1','0'),
            ('0','1','0','0','0','0','0','1','1','1','0','0','0','0'),
            ('0','1','0','0','0','0','0','1','1','1','0','0','1','0'),
            ('0','1','0','0','0','0','0','1','1','1','0','1','0','0'),
            ('0','1','0','0','0','0','0','1','1','1','0','1','1','0'),
            ('0','1','0','0','0','0','0','1','1','1','1','0','0','0'),
            ('0','1','0','0','0','0','0','1','1','1','1','0','1','0'),
            ('0','1','0','0','0','0','0','1','1','1','1','1','0','0'),
            ('0','1','0','0','0','0','0','1','1','1','1','1','1','0'),
            ('0','1','0','0','0','0','1','0','0','0','0','0','0','0'),
            ('0','1','0','0','0','0','1','0','0','0','0','0','1','0'),
            ('0','1','0','0','0','0','1','0','0','0','0','1','0','0'),
            ('0','1','0','0','0','0','1','0','0','0','0','1','1','0'),
            ('0','1','0','0','0','0','1','0','0','0','1','0','0','0'),
            ('0','1','0','0','0','0','1','0','0','0','1','0','1','0'),
            ('0','1','0','0','0','0','1','0','0','0','1','1','0','0'),
            ('0','1','0','0','0','0','1','0','0','0','1','1','1','0'),
            ('0','1','0','0','0','0','1','0','0','1','0','0','0','0'),
            ('0','1','0','0','0','0','1','0','0','1','0','0','1','0'),
            ('0','1','0','0','0','0','1','0','0','1','0','1','0','0'),
            ('0','1','0','0','0','0','1','0','0','1','0','1','1','0'),
            ('0','1','0','0','0','0','1','0','0','1','1','0','0','0'),
            ('0','1','0','0','0','0','1','0','0','1','1','0','1','0'),
            ('0','1','0','0','0','0','1','0','0','1','1','1','0','0'),
            ('0','1','0','0','0','0','1','0','0','1','1','1','1','0'),
            ('0','1','0','0','0','0','1','0','1','0','0','0','0','0'),
            ('0','1','0','0','0','0','1','0','1','0','0','0','1','0'),
            ('0','1','0','0','0','0','1','0','1','0','0','1','0','0'),
            ('0','1','0','0','0','0','1','0','1','0','0','1','1','0'),
            ('0','1','0','0','0','0','1','0','1','0','1','0','0','0'),
            ('0','1','0','0','0','0','1','0','1','0','1','0','1','0'),
            ('0','1','0','0','0','0','1','0','1','0','1','1','0','0'),
            ('0','1','0','0','0','0','1','0','1','0','1','1','1','0'),
            ('0','1','0','0','0','0','1','0','1','1','0','0','0','0'),
            ('0','1','0','0','0','0','1','0','1','1','0','0','1','0'),
            ('0','1','0','0','0','0','1','0','1','1','0','1','0','0'),
            ('0','1','0','0','0','0','1','0','1','1','0','1','1','0'),
            ('0','1','0','0','0','0','1','0','1','1','1','0','0','0'),
            ('0','1','0','0','0','0','1','0','1','1','1','0','1','0'),
            ('0','1','0','0','0','0','1','0','1','1','1','1','0','0'),
            ('0','1','0','0','0','0','1','0','1','1','1','1','1','0'),
            ('0','1','0','0','0','0','1','1','0','0','0','0','0','0'),
            ('0','1','0','0','0','0','1','1','0','0','0','0','1','0'),
            ('0','1','0','0','0','0','1','1','0','0','0','1','0','0'),
            ('0','1','0','0','0','0','1','1','0','0','0','1','1','0'),
            ('0','1','0','0','0','0','1','1','0','0','1','0','0','0'),
            ('0','1','0','0','0','0','1','1','0','0','1','0','1','0'),
            ('0','1','0','0','0','0','1','1','0','0','1','1','0','0'),
            ('0','1','0','0','0','0','1','1','0','0','1','1','1','0'),
            ('0','1','0','0','0','0','1','1','0','1','0','0','0','0'),
            ('0','1','0','0','0','0','1','1','0','1','0','0','1','0'),
            ('0','1','0','0','0','0','1','1','0','1','0','1','0','0'),
            ('0','1','0','0','0','0','1','1','0','1','0','1','1','0'),
            ('0','1','0','0','0','0','1','1','0','1','1','0','0','0'),
            ('0','1','0','0','0','0','1','1','0','1','1','0','1','0'),
            ('0','1','0','0','0','0','1','1','0','1','1','1','0','0'),
            ('0','1','0','0','0','0','1','1','0','1','1','1','1','0'),
            ('0','1','0','0','0','0','1','1','1','0','0','0','0','0'),
            ('0','1','0','0','0','0','1','1','1','0','0','0','1','0'),
            ('0','1','0','0','0','0','1','1','1','0','0','1','0','0'),
            ('0','1','0','0','0','0','1','1','1','0','0','1','1','0'),
            ('0','1','0','0','0','0','1','1','1','0','1','0','0','0'),
            ('0','1','0','0','0','0','1','1','1','0','1','0','1','0'),
            ('0','1','0','0','0','0','1','1','1','0','1','1','0','0'),
            ('0','1','0','0','0','0','1','1','1','0','1','1','1','0'),
            ('0','1','0','0','0','0','1','1','1','1','0','0','0','0'),
            ('0','1','0','0','0','0','1','1','1','1','0','0','1','0'),
            ('0','1','0','0','0','0','1','1','1','1','0','1','0','0'),
            ('0','1','0','0','0','0','1','1','1','1','0','1','1','0'),
            ('0','1','0','0','0','0','1','1','1','1','1','0','0','0'),
            ('0','1','0','0','0','0','1','1','1','1','1','0','1','0'),
            ('0','1','0','0','0','0','1','1','1','1','1','1','0','0'),
            ('0','1','0','0','0','0','1','1','1','1','1','1','1','0'),
            ('0','1','0','0','0','1','0','0','0','0','0','0','0','0'),
            ('0','1','0','0','0','1','0','0','0','0','0','0','1','0'),
            ('0','1','0','0','0','1','0','0','0','0','0','1','0','0'),
            ('0','1','0','0','0','1','0','0','0','0','0','1','1','0'),
            ('0','1','0','0','0','1','0','0','0','0','1','0','0','0'),
            ('0','1','0','0','0','1','0','0','0','0','1','0','1','0'),
            ('0','1','0','0','0','1','0','0','0','0','1','1','0','0'),
            ('0','1','0','0','0','1','0','0','0','0','1','1','1','0'),
            ('0','1','0','0','0','1','0','0','0','1','0','0','0','0'),
            ('0','1','0','0','0','1','0','0','0','1','0','0','1','0'),
            ('0','1','0','0','0','1','0','0','0','1','0','1','0','0'),
            ('0','1','0','0','0','1','0','0','0','1','0','1','1','0'),
            ('0','1','0','0','0','1','0','0','0','1','1','0','0','0'),
            ('0','1','0','0','0','1','0','0','0','1','1','0','1','0'),
            ('0','1','0','0','0','1','0','0','0','1','1','1','0','0'),
            ('0','1','0','0','0','1','0','0','0','1','1','1','1','0'),
            ('0','1','0','0','0','1','0','0','1','0','0','0','0','0'),
            ('0','1','0','0','0','1','0','0','1','0','0','0','1','0'),
            ('0','1','0','0','0','1','0','0','1','0','0','1','0','0'),
            ('0','1','0','0','0','1','0','0','1','0','0','1','1','0'),
            ('0','1','0','0','0','1','0','0','1','0','1','0','0','0'),
            ('0','1','0','0','0','1','0','0','1','0','1','0','1','0'),
            ('0','1','0','0','0','1','0','0','1','0','1','1','0','0'),
            ('0','1','0','0','0','1','0','0','1','0','1','1','1','0'),
            ('0','1','0','0','0','1','0','0','1','1','0','0','0','0'),
            ('0','1','0','0','0','1','0','0','1','1','0','0','1','0'),
            ('0','1','0','0','0','1','0','0','1','1','0','1','0','0'),
            ('0','1','0','0','0','1','0','0','1','1','0','1','1','0'),
            ('0','1','0','0','0','1','0','0','1','1','1','0','0','0'),
            ('0','1','0','0','0','1','0','0','1','1','1','0','1','0'),
            ('0','1','0','0','0','1','0','0','1','1','1','1','0','0'),
            ('0','1','0','0','0','1','0','0','1','1','1','1','1','0'),
            ('0','1','0','0','0','1','0','1','0','0','0','0','0','0'),
            ('0','1','0','0','0','1','0','1','0','0','0','0','1','0'),
            ('0','1','0','0','0','1','0','1','0','0','0','1','0','0'),
            ('0','1','0','0','0','1','0','1','0','0','0','1','1','0'),
            ('0','1','0','0','0','1','0','1','0','0','1','0','0','0'),
            ('0','1','0','0','0','1','0','1','0','0','1','0','1','0'),
            ('0','1','0','0','0','1','0','1','0','0','1','1','0','0'),
            ('0','1','0','0','0','1','0','1','0','0','1','1','1','0'),
            ('0','1','0','0','0','1','0','1','0','1','0','0','0','0'),
            ('0','1','0','0','0','1','0','1','0','1','0','0','1','0'),
            ('0','1','0','0','0','1','0','1','0','1','0','1','0','0'),
            ('0','1','0','0','0','1','0','1','0','1','0','1','1','0'),
            ('0','1','0','0','0','1','0','1','0','1','1','0','0','0'),
            ('0','1','0','0','0','1','0','1','0','1','1','0','1','0'),
            ('0','1','0','0','0','1','0','1','0','1','1','1','0','0'),
            ('0','1','0','0','0','1','0','1','0','1','1','1','1','0'),
            ('0','1','0','0','0','1','0','1','1','0','0','0','0','0'),
            ('0','1','0','0','0','1','0','1','1','0','0','0','1','0'),
            ('0','1','0','0','0','1','0','1','1','0','0','1','0','0'),
            ('0','1','0','0','0','1','0','1','1','0','0','1','1','0'),
            ('0','1','0','0','0','1','0','1','1','0','1','0','0','0'),
            ('0','1','0','0','0','1','0','1','1','0','1','0','1','0'),
            ('0','1','0','0','0','1','0','1','1','0','1','1','0','0'),
            ('0','1','0','0','0','1','0','1','1','0','1','1','1','0'),
            ('0','1','0','0','0','1','0','1','1','1','0','0','0','0'),
            ('0','1','0','0','0','1','0','1','1','1','0','0','1','0'),
            ('0','1','0','0','0','1','0','1','1','1','0','1','0','0'),
            ('0','1','0','0','0','1','0','1','1','1','0','1','1','0'),
            ('0','1','0','0','0','1','0','1','1','1','1','0','0','0'),
            ('0','1','0','0','0','1','0','1','1','1','1','0','1','0'),
            ('0','1','0','0','0','1','0','1','1','1','1','1','0','0'),
            ('0','1','0','0','0','1','0','1','1','1','1','1','1','0'),
            ('0','1','0','0','0','1','1','0','0','0','0','0','0','0'),
            ('0','1','0','0','0','1','1','0','0','0','0','0','1','0'),
            ('0','1','0','0','0','1','1','0','0','0','0','1','0','0'),
            ('0','1','0','0','0','1','1','0','0','0','0','1','1','0'),
            ('0','1','0','0','0','1','1','0','0','0','1','0','0','0'),
            ('0','1','0','0','0','1','1','0','0','0','1','0','1','0'),
            ('0','1','0','0','0','1','1','0','0','0','1','1','0','0'),
            ('0','1','0','0','0','1','1','0','0','0','1','1','1','0'),
            ('0','1','0','0','0','1','1','0','0','1','0','0','0','0'),
            ('0','1','0','0','0','1','1','0','0','1','0','0','1','0'),
            ('0','1','0','0','0','1','1','0','0','1','0','1','0','0'),
            ('0','1','0','0','0','1','1','0','0','1','0','1','1','0'),
            ('0','1','0','0','0','1','1','0','0','1','1','0','0','0'),
            ('0','1','0','0','0','1','1','0','0','1','1','0','1','0'),
            ('0','1','0','0','0','1','1','0','0','1','1','1','0','0'),
            ('0','1','0','0','0','1','1','0','0','1','1','1','1','0'),
            ('0','1','0','0','0','1','1','0','1','0','0','0','0','0'),
            ('0','1','0','0','0','1','1','0','1','0','0','0','1','0'),
            ('0','1','0','0','0','1','1','0','1','0','0','1','0','0'),
            ('0','1','0','0','0','1','1','0','1','0','0','1','1','0'),
            ('0','1','0','0','0','1','1','0','1','0','1','0','0','0'),
            ('0','1','0','0','0','1','1','0','1','0','1','0','1','0'),
            ('0','1','0','0','0','1','1','0','1','0','1','1','0','0'),
            ('0','1','0','0','0','1','1','0','1','0','1','1','1','0'),
            ('0','1','0','0','0','1','1','0','1','1','0','0','0','0'),
            ('0','1','0','0','0','1','1','0','1','1','0','0','1','0'),
            ('0','1','0','0','0','1','1','0','1','1','0','1','0','0'),
            ('0','1','0','0','0','1','1','0','1','1','0','1','1','0'),
            ('0','1','0','0','0','1','1','0','1','1','1','0','0','0'),
            ('0','1','0','0','0','1','1','0','1','1','1','0','1','0'),
            ('0','1','0','0','0','1','1','0','1','1','1','1','0','0'),
            ('0','1','0','0','0','1','1','0','1','1','1','1','1','0'),
            ('0','1','0','0','0','1','1','1','0','0','0','0','0','0'),
            ('0','1','0','0','0','1','1','1','0','0','0','0','1','0'),
            ('0','1','0','0','0','1','1','1','0','0','0','1','0','0'),
            ('0','1','0','0','0','1','1','1','0','0','0','1','1','0'),
            ('0','1','0','0','0','1','1','1','0','0','1','0','0','0'),
            ('0','1','0','0','0','1','1','1','0','0','1','0','1','0'),
            ('0','1','0','0','0','1','1','1','0','0','1','1','0','0'),
            ('0','1','0','0','0','1','1','1','0','0','1','1','1','0'),
            ('0','1','0','0','0','1','1','1','0','1','0','0','0','0'),
            ('0','1','0','0','0','1','1','1','0','1','0','0','1','0'),
            ('0','1','0','0','0','1','1','1','0','1','0','1','0','0'),
            ('0','1','0','0','0','1','1','1','0','1','0','1','1','0'),
            ('0','1','0','0','0','1','1','1','0','1','1','0','0','0'),
            ('0','1','0','0','0','1','1','1','0','1','1','0','1','0'),
            ('0','1','0','0','0','1','1','1','0','1','1','1','0','0'),
            ('0','1','0','0','0','1','1','1','0','1','1','1','1','0'),
            ('0','1','0','0','0','1','1','1','1','0','0','0','0','0'),
            ('0','1','0','0','0','1','1','1','1','0','0','0','1','0'),
            ('0','1','0','0','0','1','1','1','1','0','0','1','0','0'),
            ('0','1','0','0','0','1','1','1','1','0','0','1','1','0'),
            ('0','1','0','0','0','1','1','1','1','0','1','0','0','0'),
            ('0','1','0','0','0','1','1','1','1','0','1','0','1','0'),
            ('0','1','0','0','0','1','1','1','1','0','1','1','0','0'),
            ('0','1','0','0','0','1','1','1','1','0','1','1','1','0'),
            ('0','1','0','0','0','1','1','1','1','1','0','0','0','0'),
            ('0','1','0','0','0','1','1','1','1','1','0','0','1','0'),
            ('0','1','0','0','0','1','1','1','1','1','0','1','0','0'),
            ('0','1','0','0','0','1','1','1','1','1','0','1','1','0'),
            ('0','1','0','0','0','1','1','1','1','1','1','0','0','0'),
            ('0','1','0','0','0','1','1','1','1','1','1','0','1','0'),
            ('0','1','0','0','0','1','1','1','1','1','1','1','0','0'),
            ('0','1','0','0','0','1','1','1','1','1','1','1','1','0'),
            ('0','1','0','0','1','0','0','0','0','0','0','0','0','0'),
            ('0','1','0','0','1','0','0','0','0','0','0','0','1','0'),
            ('0','1','0','0','1','0','0','0','0','0','0','1','0','0'),
            ('0','1','0','0','1','0','0','0','0','0','0','1','1','0'),
            ('0','1','0','0','1','0','0','0','0','0','1','0','0','0'),
            ('0','1','0','0','1','0','0','0','0','0','1','0','1','0'),
            ('0','1','0','0','1','0','0','0','0','0','1','1','0','0'),
            ('0','1','0','0','1','0','0','0','0','0','1','1','1','0'),
            ('0','1','0','0','1','0','0','0','0','1','0','0','0','0'),
            ('0','1','0','0','1','0','0','0','0','1','0','0','1','0'),
            ('0','1','0','0','1','0','0','0','0','1','0','1','0','0'),
            ('0','1','0','0','1','0','0','0','0','1','0','1','1','0'),
            ('0','1','0','0','1','0','0','0','0','1','1','0','0','0'),
            ('0','1','0','0','1','0','0','0','0','1','1','0','1','0'),
            ('0','1','0','0','1','0','0','0','0','1','1','1','0','0'),
            ('0','1','0','0','1','0','0','0','0','1','1','1','1','0'),
            ('0','1','0','0','1','0','0','0','1','0','0','0','0','0'),
            ('0','1','0','0','1','0','0','0','1','0','0','0','1','0'),
            ('0','1','0','0','1','0','0','0','1','0','0','1','0','0'),
            ('0','1','0','0','1','0','0','0','1','0','0','1','1','0'),
            ('0','1','0','0','1','0','0','0','1','0','1','0','0','0'),
            ('0','1','0','0','1','0','0','0','1','0','1','0','1','0'),
            ('0','1','0','0','1','0','0','0','1','0','1','1','0','0'),
            ('0','1','0','0','1','0','0','0','1','0','1','1','1','0'),
            ('0','1','0','0','1','0','0','0','1','1','0','0','0','0'),
            ('0','1','0','0','1','0','0','0','1','1','0','0','1','0'),
            ('0','1','0','0','1','0','0','0','1','1','0','1','0','0'),
            ('0','1','0','0','1','0','0','0','1','1','0','1','1','0'),
            ('0','1','0','0','1','0','0','0','1','1','1','0','0','0'),
            ('0','1','0','0','1','0','0','0','1','1','1','0','1','0'),
            ('0','1','0','0','1','0','0','0','1','1','1','1','0','0'),
            ('0','1','0','0','1','0','0','0','1','1','1','1','1','0'),
            ('0','1','0','0','1','0','0','1','0','0','0','0','0','0'),
            ('0','1','0','0','1','0','0','1','0','0','0','0','1','0'),
            ('0','1','0','0','1','0','0','1','0','0','0','1','0','0'),
            ('0','1','0','0','1','0','0','1','0','0','0','1','1','0'),
            ('0','1','0','0','1','0','0','1','0','0','1','0','0','0'),
            ('0','1','0','0','1','0','0','1','0','0','1','0','1','0'),
            ('0','1','0','0','1','0','0','1','0','0','1','1','0','0'),
            ('0','1','0','0','1','0','0','1','0','0','1','1','1','0'),
            ('0','1','0','0','1','0','0','1','0','1','0','0','0','0'),
            ('0','1','0','0','1','0','0','1','0','1','0','0','1','0'),
            ('0','1','0','0','1','0','0','1','0','1','0','1','0','0'),
            ('0','1','0','0','1','0','0','1','0','1','0','1','1','0'),
            ('0','1','0','0','1','0','0','1','0','1','1','0','0','0'),
            ('0','1','0','0','1','0','0','1','0','1','1','0','1','0'),
            ('0','1','0','0','1','0','0','1','0','1','1','1','0','0'),
            ('0','1','0','0','1','0','0','1','0','1','1','1','1','0'),
            ('0','1','0','0','1','0','0','1','1','0','0','0','0','0'),
            ('0','1','0','0','1','0','0','1','1','0','0','0','1','0'),
            ('0','1','0','0','1','0','0','1','1','0','0','1','0','0'),
            ('0','1','0','0','1','0','0','1','1','0','0','1','1','0'),
            ('0','1','0','0','1','0','0','1','1','0','1','0','0','0'),
            ('0','1','0','0','1','0','0','1','1','0','1','0','1','0'),
            ('0','1','0','0','1','0','0','1','1','0','1','1','0','0'),
            ('0','1','0','0','1','0','0','1','1','0','1','1','1','0'),
            ('0','1','0','0','1','0','0','1','1','1','0','0','0','0'),
            ('0','1','0','0','1','0','0','1','1','1','0','0','1','0'),
            ('0','1','0','0','1','0','0','1','1','1','0','1','0','0'),
            ('0','1','0','0','1','0','0','1','1','1','0','1','1','0'),
            ('0','1','0','0','1','0','0','1','1','1','1','0','0','0'),
            ('0','1','0','0','1','0','0','1','1','1','1','0','1','0'),
            ('0','1','0','0','1','0','0','1','1','1','1','1','0','0'),
            ('0','1','0','0','1','0','0','1','1','1','1','1','1','0'),
            ('0','1','0','0','1','0','1','0','0','0','0','0','0','0'),
            ('0','1','0','0','1','0','1','0','0','0','0','0','1','0'),
            ('0','1','0','0','1','0','1','0','0','0','0','1','0','0'),
            ('0','1','0','0','1','0','1','0','0','0','0','1','1','0'),
            ('0','1','0','0','1','0','1','0','0','0','1','0','0','0'),
            ('0','1','0','0','1','0','1','0','0','0','1','0','1','0'),
            ('0','1','0','0','1','0','1','0','0','0','1','1','0','0'),
            ('0','1','0','0','1','0','1','0','0','0','1','1','1','0'),
            ('0','1','0','0','1','0','1','0','0','1','0','0','0','0'),
            ('0','1','0','0','1','0','1','0','0','1','0','0','1','0'),
            ('0','1','0','0','1','0','1','0','0','1','0','1','0','0'),
            ('0','1','0','0','1','0','1','0','0','1','0','1','1','0'),
            ('0','1','0','0','1','0','1','0','0','1','1','0','0','0'),
            ('0','1','0','0','1','0','1','0','0','1','1','0','1','0'),
            ('0','1','0','0','1','0','1','0','0','1','1','1','0','0'),
            ('0','1','0','0','1','0','1','0','0','1','1','1','1','0'),
            ('0','1','0','0','1','0','1','0','1','0','0','0','0','0'),
            ('0','1','0','0','1','0','1','0','1','0','0','0','1','0'),
            ('0','1','0','0','1','0','1','0','1','0','0','1','0','0'),
            ('0','1','0','0','1','0','1','0','1','0','0','1','1','0'),
            ('0','1','0','0','1','0','1','0','1','0','1','0','0','0'),
            ('0','1','0','0','1','0','1','0','1','0','1','0','1','0'),
            ('0','1','0','0','1','0','1','0','1','0','1','1','0','0'),
            ('0','1','0','0','1','0','1','0','1','0','1','1','1','0'),
            ('0','1','0','0','1','0','1','0','1','1','0','0','0','0'),
            ('0','1','0','0','1','0','1','0','1','1','0','0','1','0'),
            ('0','1','0','0','1','0','1','0','1','1','0','1','0','0'),
            ('0','1','0','0','1','0','1','0','1','1','0','1','1','0'),
            ('0','1','0','0','1','0','1','0','1','1','1','0','0','0'),
            ('0','1','0','0','1','0','1','0','1','1','1','0','1','0'),
            ('0','1','0','0','1','0','1','0','1','1','1','1','0','0'),
            ('0','1','0','0','1','0','1','0','1','1','1','1','1','0'),
            ('0','1','0','0','1','0','1','1','0','0','0','0','0','0'),
            ('0','1','0','0','1','0','1','1','0','0','0','0','1','0'),
            ('0','1','0','0','1','0','1','1','0','0','0','1','0','0'),
            ('0','1','0','0','1','0','1','1','0','0','0','1','1','0'),
            ('0','1','0','0','1','0','1','1','0','0','1','0','0','0'),
            ('0','1','0','0','1','0','1','1','0','0','1','0','1','0'),
            ('0','1','0','0','1','0','1','1','0','0','1','1','0','0'),
            ('0','1','0','0','1','0','1','1','0','0','1','1','1','0'),
            ('0','1','0','0','1','0','1','1','0','1','0','0','0','0'),
            ('0','1','0','0','1','0','1','1','0','1','0','0','1','0'),
            ('0','1','0','0','1','0','1','1','0','1','0','1','0','0'),
            ('0','1','0','0','1','0','1','1','0','1','0','1','1','0'),
            ('0','1','0','0','1','0','1','1','0','1','1','0','0','0'),
            ('0','1','0','0','1','0','1','1','0','1','1','0','1','0'),
            ('0','1','0','0','1','0','1','1','0','1','1','1','0','0'),
            ('0','1','0','0','1','0','1','1','0','1','1','1','1','0'),
            ('0','1','0','0','1','0','1','1','1','0','0','0','0','0'),
            ('0','1','0','0','1','0','1','1','1','0','0','0','1','0'),
            ('0','1','0','0','1','0','1','1','1','0','0','1','0','0'),
            ('0','1','0','0','1','0','1','1','1','0','0','1','1','0'),
            ('0','1','0','0','1','0','1','1','1','0','1','0','0','0'),
            ('0','1','0','0','1','0','1','1','1','0','1','0','1','0'),
            ('0','1','0','0','1','0','1','1','1','0','1','1','0','0'),
            ('0','1','0','0','1','0','1','1','1','0','1','1','1','0'),
            ('0','1','0','0','1','0','1','1','1','1','0','0','0','0'),
            ('0','1','0','0','1','0','1','1','1','1','0','0','1','0'),
            ('0','1','0','0','1','0','1','1','1','1','0','1','0','0'),
            ('0','1','0','0','1','0','1','1','1','1','0','1','1','0'),
            ('0','1','0','0','1','0','1','1','1','1','1','0','0','0'),
            ('0','1','0','0','1','0','1','1','1','1','1','0','1','0'),
            ('0','1','0','0','1','0','1','1','1','1','1','1','0','0'),
            ('0','1','0','0','1','0','1','1','1','1','1','1','1','0'),
            ('0','1','0','0','1','1','0','0','0','0','0','0','0','0'),
            ('0','1','0','0','1','1','0','0','0','0','0','0','1','0'),
            ('0','1','0','0','1','1','0','0','0','0','0','1','0','0'),
            ('0','1','0','0','1','1','0','0','0','0','0','1','1','0'),
            ('0','1','0','0','1','1','0','0','0','0','1','0','0','0'),
            ('0','1','0','0','1','1','0','0','0','0','1','0','1','0'),
            ('0','1','0','0','1','1','0','0','0','0','1','1','0','0'),
            ('0','1','0','0','1','1','0','0','0','0','1','1','1','0'),
            ('0','1','0','0','1','1','0','0','0','1','0','0','0','0'),
            ('0','1','0','0','1','1','0','0','0','1','0','0','1','0'),
            ('0','1','0','0','1','1','0','0','0','1','0','1','0','0'),
            ('0','1','0','0','1','1','0','0','0','1','0','1','1','0'),
            ('0','1','0','0','1','1','0','0','0','1','1','0','0','0'),
            ('0','1','0','0','1','1','0','0','0','1','1','0','1','0'),
            ('0','1','0','0','1','1','0','0','0','1','1','1','0','0'),
            ('0','1','0','0','1','1','0','0','0','1','1','1','1','0'),
            ('0','1','0','0','1','1','0','0','1','0','0','0','0','0'),
            ('0','1','0','0','1','1','0','0','1','0','0','0','1','0'),
            ('0','1','0','0','1','1','0','0','1','0','0','1','0','0'),
            ('0','1','0','0','1','1','0','0','1','0','0','1','1','0'),
            ('0','1','0','0','1','1','0','0','1','0','1','0','0','0'),
            ('0','1','0','0','1','1','0','0','1','0','1','0','1','0'),
            ('0','1','0','0','1','1','0','0','1','0','1','1','0','0'),
            ('0','1','0','0','1','1','0','0','1','0','1','1','1','0'),
            ('0','1','0','0','1','1','0','0','1','1','0','0','0','0'),
            ('0','1','0','0','1','1','0','0','1','1','0','0','1','0'),
            ('0','1','0','0','1','1','0','0','1','1','0','1','0','0'),
            ('0','1','0','0','1','1','0','0','1','1','0','1','1','0'),
            ('0','1','0','0','1','1','0','0','1','1','1','0','0','0'),
            ('0','1','0','0','1','1','0','0','1','1','1','0','1','0'),
            ('0','1','0','0','1','1','0','0','1','1','1','1','0','0'),
            ('0','1','0','0','1','1','0','0','1','1','1','1','1','0'),
            ('0','1','0','0','1','1','0','1','0','0','0','0','0','0'),
            ('0','1','0','0','1','1','0','1','0','0','0','0','1','0'),
            ('0','1','0','0','1','1','0','1','0','0','0','1','0','0'),
            ('0','1','0','0','1','1','0','1','0','0','0','1','1','0'),
            ('0','1','0','0','1','1','0','1','0','0','1','0','0','0'),
            ('0','1','0','0','1','1','0','1','0','0','1','0','1','0'),
            ('0','1','0','0','1','1','0','1','0','0','1','1','0','0'),
            ('0','1','0','0','1','1','0','1','0','0','1','1','1','0'),
            ('0','1','0','0','1','1','0','1','0','1','0','0','0','0'),
            ('0','1','0','0','1','1','0','1','0','1','0','0','1','0'),
            ('0','1','0','0','1','1','0','1','0','1','0','1','0','0'),
            ('0','1','0','0','1','1','0','1','0','1','0','1','1','0'),
            ('0','1','0','0','1','1','0','1','0','1','1','0','0','0'),
            ('0','1','0','0','1','1','0','1','0','1','1','0','1','0'),
            ('0','1','0','0','1','1','0','1','0','1','1','1','0','0'),
            ('0','1','0','0','1','1','0','1','0','1','1','1','1','0'),
            ('0','1','0','0','1','1','0','1','1','0','0','0','0','0'),
            ('0','1','0','0','1','1','0','1','1','0','0','0','1','0'),
            ('0','1','0','0','1','1','0','1','1','0','0','1','0','0'),
            ('0','1','0','0','1','1','0','1','1','0','0','1','1','0'),
            ('0','1','0','0','1','1','0','1','1','0','1','0','0','0'),
            ('0','1','0','0','1','1','0','1','1','0','1','0','1','0'),
            ('0','1','0','0','1','1','0','1','1','0','1','1','0','0'),
            ('0','1','0','0','1','1','0','1','1','0','1','1','1','0'),
            ('0','1','0','0','1','1','0','1','1','1','0','0','0','0'),
            ('0','1','0','0','1','1','0','1','1','1','0','0','1','0'),
            ('0','1','0','0','1','1','0','1','1','1','0','1','0','0'),
            ('0','1','0','0','1','1','0','1','1','1','0','1','1','0'),
            ('0','1','0','0','1','1','0','1','1','1','1','0','0','0'),
            ('0','1','0','0','1','1','0','1','1','1','1','0','1','0'),
            ('0','1','0','0','1','1','0','1','1','1','1','1','0','0'),
            ('0','1','0','0','1','1','0','1','1','1','1','1','1','0'),
            ('0','1','0','0','1','1','1','0','0','0','0','0','0','0'),
            ('0','1','0','0','1','1','1','0','0','0','0','0','1','0'),
            ('0','1','0','0','1','1','1','0','0','0','0','1','0','0'),
            ('0','1','0','0','1','1','1','0','0','0','0','1','1','0'),
            ('0','1','0','0','1','1','1','0','0','0','1','0','0','0'),
            ('0','1','0','0','1','1','1','0','0','0','1','0','1','0'),
            ('0','1','0','0','1','1','1','0','0','0','1','1','0','0'),
            ('0','1','0','0','1','1','1','0','0','0','1','1','1','0'),
            ('0','1','0','0','1','1','1','0','0','1','0','0','0','0'),
            ('0','1','0','0','1','1','1','0','0','1','0','0','1','0'),
            ('0','1','0','0','1','1','1','0','0','1','0','1','0','0'),
            ('0','1','0','0','1','1','1','0','0','1','0','1','1','0'),
            ('0','1','0','0','1','1','1','0','0','1','1','0','0','0'),
            ('0','1','0','0','1','1','1','0','0','1','1','0','1','0'),
            ('0','1','0','0','1','1','1','0','0','1','1','1','0','0'),
            ('0','1','0','0','1','1','1','0','0','1','1','1','1','0'),
            ('0','1','0','0','1','1','1','0','1','0','0','0','0','0'),
            ('0','1','0','0','1','1','1','0','1','0','0','0','1','0'),
            ('0','1','0','0','1','1','1','0','1','0','0','1','0','0'),
            ('0','1','0','0','1','1','1','0','1','0','0','1','1','0'),
            ('0','1','0','0','1','1','1','0','1','0','1','0','0','0'),
            ('0','1','0','0','1','1','1','0','1','0','1','0','1','0'),
            ('0','1','0','0','1','1','1','0','1','0','1','1','0','0'),
            ('0','1','0','0','1','1','1','0','1','0','1','1','1','0'),
            ('0','1','0','0','1','1','1','0','1','1','0','0','0','0'),
            ('0','1','0','0','1','1','1','0','1','1','0','0','1','0'),
            ('0','1','0','0','1','1','1','0','1','1','0','1','0','0'),
            ('0','1','0','0','1','1','1','0','1','1','0','1','1','0'),
            ('0','1','0','0','1','1','1','0','1','1','1','0','0','0'),
            ('0','1','0','0','1','1','1','0','1','1','1','0','1','0'),
            ('0','1','0','0','1','1','1','0','1','1','1','1','0','0'),
            ('0','1','0','0','1','1','1','0','1','1','1','1','1','0'),
            ('0','1','0','0','1','1','1','1','0','0','0','0','0','0'),
            ('0','1','0','0','1','1','1','1','0','0','0','0','1','0'),
            ('0','1','0','0','1','1','1','1','0','0','0','1','0','0'),
            ('0','1','0','0','1','1','1','1','0','0','0','1','1','0'),
            ('0','1','0','0','1','1','1','1','0','0','1','0','0','0'),
            ('0','1','0','0','1','1','1','1','0','0','1','0','1','0'),
            ('0','1','0','0','1','1','1','1','0','0','1','1','0','0'),
            ('0','1','0','0','1','1','1','1','0','0','1','1','1','0'),
            ('0','1','0','0','1','1','1','1','0','1','0','0','0','0'),
            ('0','1','0','0','1','1','1','1','0','1','0','0','1','0'),
            ('0','1','0','0','1','1','1','1','0','1','0','1','0','0'),
            ('0','1','0','0','1','1','1','1','0','1','0','1','1','0'),
            ('0','1','0','0','1','1','1','1','0','1','1','0','0','0'),
            ('0','1','0','0','1','1','1','1','0','1','1','0','1','0'),
            ('0','1','0','0','1','1','1','1','0','1','1','1','0','0'),
            ('0','1','0','0','1','1','1','1','0','1','1','1','1','0'),
            ('0','1','0','0','1','1','1','1','1','0','0','0','0','0'),
            ('0','1','0','0','1','1','1','1','1','0','0','0','1','0'),
            ('0','1','0','0','1','1','1','1','1','0','0','1','0','0'),
            ('0','1','0','0','1','1','1','1','1','0','0','1','1','0'),
            ('0','1','0','0','1','1','1','1','1','0','1','0','0','0'),
            ('0','1','0','0','1','1','1','1','1','0','1','0','1','0'),
            ('0','1','0','0','1','1','1','1','1','0','1','1','0','0'),
            ('0','1','0','0','1','1','1','1','1','0','1','1','1','0'),
            ('0','1','0','0','1','1','1','1','1','1','0','0','0','0'),
            ('0','1','0','0','1','1','1','1','1','1','0','0','1','0'),
            ('0','1','0','0','1','1','1','1','1','1','0','1','0','0'),
            ('0','1','0','0','1','1','1','1','1','1','0','1','1','0'),
            ('0','1','0','0','1','1','1','1','1','1','1','0','0','0'),
            ('0','1','0','0','1','1','1','1','1','1','1','0','1','0'),
            ('0','1','0','0','1','1','1','1','1','1','1','1','0','0'),
            ('0','1','0','0','1','1','1','1','1','1','1','1','1','0'),
            ('0','1','0','1','0','0','0','0','0','0','0','0','0','0'),
            ('0','1','0','1','0','0','0','0','0','0','0','0','1','0'),
            ('0','1','0','1','0','0','0','0','0','0','0','1','0','0'),
            ('0','1','0','1','0','0','0','0','0','0','0','1','1','0'),
            ('0','1','0','1','0','0','0','0','0','0','1','0','0','0'),
            ('0','1','0','1','0','0','0','0','0','0','1','0','1','0'),
            ('0','1','0','1','0','0','0','0','0','0','1','1','0','0'),
            ('0','1','0','1','0','0','0','0','0','0','1','1','1','0'),
            ('0','1','0','1','0','0','0','0','0','1','0','0','0','0'),
            ('0','1','0','1','0','0','0','0','0','1','0','0','1','0'),
            ('0','1','0','1','0','0','0','0','0','1','0','1','0','0'),
            ('0','1','0','1','0','0','0','0','0','1','0','1','1','0'),
            ('0','1','0','1','0','0','0','0','0','1','1','0','0','0'),
            ('0','1','0','1','0','0','0','0','0','1','1','0','1','0'),
            ('0','1','0','1','0','0','0','0','0','1','1','1','0','0'),
            ('0','1','0','1','0','0','0','0','0','1','1','1','1','0'),
            ('0','1','0','1','0','0','0','0','1','0','0','0','0','0'),
            ('0','1','0','1','0','0','0','0','1','0','0','0','1','0'),
            ('0','1','0','1','0','0','0','0','1','0','0','1','0','0'),
            ('0','1','0','1','0','0','0','0','1','0','0','1','1','0'),
            ('0','1','0','1','0','0','0','0','1','0','1','0','0','0'),
            ('0','1','0','1','0','0','0','0','1','0','1','0','1','0'),
            ('0','1','0','1','0','0','0','0','1','0','1','1','0','0'),
            ('0','1','0','1','0','0','0','0','1','0','1','1','1','0'),
            ('0','1','0','1','0','0','0','0','1','1','0','0','0','0'),
            ('0','1','0','1','0','0','0','0','1','1','0','0','1','0'),
            ('0','1','0','1','0','0','0','0','1','1','0','1','0','0'),
            ('0','1','0','1','0','0','0','0','1','1','0','1','1','0'),
            ('0','1','0','1','0','0','0','0','1','1','1','0','0','0'),
            ('0','1','0','1','0','0','0','0','1','1','1','0','1','0'),
            ('0','1','0','1','0','0','0','0','1','1','1','1','0','0'),
            ('0','1','0','1','0','0','0','0','1','1','1','1','1','0'),
            ('0','1','0','1','0','0','0','1','0','0','0','0','0','0'),
            ('0','1','0','1','0','0','0','1','0','0','0','0','1','0'),
            ('0','1','0','1','0','0','0','1','0','0','0','1','0','0'),
            ('0','1','0','1','0','0','0','1','0','0','0','1','1','0'),
            ('0','1','0','1','0','0','0','1','0','0','1','0','0','0'),
            ('0','1','0','1','0','0','0','1','0','0','1','0','1','0'),
            ('0','1','0','1','0','0','0','1','0','0','1','1','0','0'),
            ('0','1','0','1','0','0','0','1','0','0','1','1','1','0'),
            ('0','1','0','1','0','0','0','1','0','1','0','0','0','0'),
            ('0','1','0','1','0','0','0','1','0','1','0','0','1','0'),
            ('0','1','0','1','0','0','0','1','0','1','0','1','0','0'),
            ('0','1','0','1','0','0','0','1','0','1','0','1','1','0'),
            ('0','1','0','1','0','0','0','1','0','1','1','0','0','0'),
            ('0','1','0','1','0','0','0','1','0','1','1','0','1','0'),
            ('0','1','0','1','0','0','0','1','0','1','1','1','0','0'),
            ('0','1','0','1','0','0','0','1','0','1','1','1','1','0'),
            ('0','1','0','1','0','0','0','1','1','0','0','0','0','0'),
            ('0','1','0','1','0','0','0','1','1','0','0','0','1','0'),
            ('0','1','0','1','0','0','0','1','1','0','0','1','0','0'),
            ('0','1','0','1','0','0','0','1','1','0','0','1','1','0'),
            ('0','1','0','1','0','0','0','1','1','0','1','0','0','0'),
            ('0','1','0','1','0','0','0','1','1','0','1','0','1','0'),
            ('0','1','0','1','0','0','0','1','1','0','1','1','0','0'),
            ('0','1','0','1','0','0','0','1','1','0','1','1','1','0'),
            ('0','1','0','1','0','0','0','1','1','1','0','0','0','0'),
            ('0','1','0','1','0','0','0','1','1','1','0','0','1','0'),
            ('0','1','0','1','0','0','0','1','1','1','0','1','0','0'),
            ('0','1','0','1','0','0','0','1','1','1','0','1','1','0'),
            ('0','1','0','1','0','0','0','1','1','1','1','0','0','0'),
            ('0','1','0','1','0','0','0','1','1','1','1','0','1','0'),
            ('0','1','0','1','0','0','0','1','1','1','1','1','0','0'),
            ('0','1','0','1','0','0','0','1','1','1','1','1','1','0'),
            ('0','1','0','1','0','0','1','0','0','0','0','0','0','0'),
            ('0','1','0','1','0','0','1','0','0','0','0','0','1','0'),
            ('0','1','0','1','0','0','1','0','0','0','0','1','0','0'),
            ('0','1','0','1','0','0','1','0','0','0','0','1','1','0'),
            ('0','1','0','1','0','0','1','0','0','0','1','0','0','0'),
            ('0','1','0','1','0','0','1','0','0','0','1','0','1','0'),
            ('0','1','0','1','0','0','1','0','0','0','1','1','0','0'),
            ('0','1','0','1','0','0','1','0','0','0','1','1','1','0'),
            ('0','1','0','1','0','0','1','0','0','1','0','0','0','0'),
            ('0','1','0','1','0','0','1','0','0','1','0','0','1','0'),
            ('0','1','0','1','0','0','1','0','0','1','0','1','0','0'),
            ('0','1','0','1','0','0','1','0','0','1','0','1','1','0'),
            ('0','1','0','1','0','0','1','0','0','1','1','0','0','0'),
            ('0','1','0','1','0','0','1','0','0','1','1','0','1','0'),
            ('0','1','0','1','0','0','1','0','0','1','1','1','0','0'),
            ('0','1','0','1','0','0','1','0','0','1','1','1','1','0'),
            ('0','1','0','1','0','0','1','0','1','0','0','0','0','0'),
            ('0','1','0','1','0','0','1','0','1','0','0','0','1','0'),
            ('0','1','0','1','0','0','1','0','1','0','0','1','0','0'),
            ('0','1','0','1','0','0','1','0','1','0','0','1','1','0'),
            ('0','1','0','1','0','0','1','0','1','0','1','0','0','0'),
            ('0','1','0','1','0','0','1','0','1','0','1','0','1','0'),
            ('0','1','0','1','0','0','1','0','1','0','1','1','0','0'),
            ('0','1','0','1','0','0','1','0','1','0','1','1','1','0'),
            ('0','1','0','1','0','0','1','0','1','1','0','0','0','0'),
            ('0','1','0','1','0','0','1','0','1','1','0','0','1','0'),
            ('0','1','0','1','0','0','1','0','1','1','0','1','0','0'),
            ('0','1','0','1','0','0','1','0','1','1','0','1','1','0'),
            ('0','1','0','1','0','0','1','0','1','1','1','0','0','0'),
            ('0','1','0','1','0','0','1','0','1','1','1','0','1','0'),
            ('0','1','0','1','0','0','1','0','1','1','1','1','0','0'),
            ('0','1','0','1','0','0','1','0','1','1','1','1','1','0'),
            ('0','1','0','1','0','0','1','1','0','0','0','0','0','0'),
            ('0','1','0','1','0','0','1','1','0','0','0','0','1','0'),
            ('0','1','0','1','0','0','1','1','0','0','0','1','0','0'),
            ('0','1','0','1','0','0','1','1','0','0','0','1','1','0'),
            ('0','1','0','1','0','0','1','1','0','0','1','0','0','0'),
            ('0','1','0','1','0','0','1','1','0','0','1','0','1','0'),
            ('0','1','0','1','0','0','1','1','0','0','1','1','0','0'),
            ('0','1','0','1','0','0','1','1','0','0','1','1','1','0'),
            ('0','1','0','1','0','0','1','1','0','1','0','0','0','0'),
            ('0','1','0','1','0','0','1','1','0','1','0','0','1','0'),
            ('0','1','0','1','0','0','1','1','0','1','0','1','0','0'),
            ('0','1','0','1','0','0','1','1','0','1','0','1','1','0'),
            ('0','1','0','1','0','0','1','1','0','1','1','0','0','0'),
            ('0','1','0','1','0','0','1','1','0','1','1','0','1','0'),
            ('0','1','0','1','0','0','1','1','0','1','1','1','0','0'),
            ('0','1','0','1','0','0','1','1','0','1','1','1','1','0'),
            ('0','1','0','1','0','0','1','1','1','0','0','0','0','0'),
            ('0','1','0','1','0','0','1','1','1','0','0','0','1','0'),
            ('0','1','0','1','0','0','1','1','1','0','0','1','0','0'),
            ('0','1','0','1','0','0','1','1','1','0','0','1','1','0'),
            ('0','1','0','1','0','0','1','1','1','0','1','0','0','0'),
            ('0','1','0','1','0','0','1','1','1','0','1','0','1','0'),
            ('0','1','0','1','0','0','1','1','1','0','1','1','0','0'),
            ('0','1','0','1','0','0','1','1','1','0','1','1','1','0'),
            ('0','1','0','1','0','0','1','1','1','1','0','0','0','0'),
            ('0','1','0','1','0','0','1','1','1','1','0','0','1','0'),
            ('0','1','0','1','0','0','1','1','1','1','0','1','0','0'),
            ('0','1','0','1','0','0','1','1','1','1','0','1','1','0'),
            ('0','1','0','1','0','0','1','1','1','1','1','0','0','0'),
            ('0','1','0','1','0','0','1','1','1','1','1','0','1','0'),
            ('0','1','0','1','0','0','1','1','1','1','1','1','0','0'),
            ('0','1','0','1','0','0','1','1','1','1','1','1','1','0'),
            ('0','1','0','1','0','1','0','0','0','0','0','0','0','0'),
            ('0','1','0','1','0','1','0','0','0','0','0','0','1','0'),
            ('0','1','0','1','0','1','0','0','0','0','0','1','0','0'),
            ('0','1','0','1','0','1','0','0','0','0','0','1','1','0'),
            ('0','1','0','1','0','1','0','0','0','0','1','0','0','0'),
            ('0','1','0','1','0','1','0','0','0','0','1','0','1','0'),
            ('0','1','0','1','0','1','0','0','0','0','1','1','0','0'),
            ('0','1','0','1','0','1','0','0','0','0','1','1','1','0'),
            ('0','1','0','1','0','1','0','0','0','1','0','0','0','0'),
            ('0','1','0','1','0','1','0','0','0','1','0','0','1','0'),
            ('0','1','0','1','0','1','0','0','0','1','0','1','0','0'),
            ('0','1','0','1','0','1','0','0','0','1','0','1','1','0'),
            ('0','1','0','1','0','1','0','0','0','1','1','0','0','0'),
            ('0','1','0','1','0','1','0','0','0','1','1','0','1','0'),
            ('0','1','0','1','0','1','0','0','0','1','1','1','0','0'),
            ('0','1','0','1','0','1','0','0','0','1','1','1','1','0'),
            ('0','1','0','1','0','1','0','0','1','0','0','0','0','0'),
            ('0','1','0','1','0','1','0','0','1','0','0','0','1','0'),
            ('0','1','0','1','0','1','0','0','1','0','0','1','0','0'),
            ('0','1','0','1','0','1','0','0','1','0','0','1','1','0'),
            ('0','1','0','1','0','1','0','0','1','0','1','0','0','0'),
            ('0','1','0','1','0','1','0','0','1','0','1','0','1','0'),
            ('0','1','0','1','0','1','0','0','1','0','1','1','0','0'),
            ('0','1','0','1','0','1','0','0','1','0','1','1','1','0'),
            ('0','1','0','1','0','1','0','0','1','1','0','0','0','0'),
            ('0','1','0','1','0','1','0','0','1','1','0','0','1','0'),
            ('0','1','0','1','0','1','0','0','1','1','0','1','0','0'),
            ('0','1','0','1','0','1','0','0','1','1','0','1','1','0'),
            ('0','1','0','1','0','1','0','0','1','1','1','0','0','0'),
            ('0','1','0','1','0','1','0','0','1','1','1','0','1','0'),
            ('0','1','0','1','0','1','0','0','1','1','1','1','0','0'),
            ('0','1','0','1','0','1','0','0','1','1','1','1','1','0'),
            ('0','1','0','1','0','1','0','1','0','0','0','0','0','0'),
            ('0','1','0','1','0','1','0','1','0','0','0','0','1','0'),
            ('0','1','0','1','0','1','0','1','0','0','0','1','0','0'),
            ('0','1','0','1','0','1','0','1','0','0','0','1','1','0'),
            ('0','1','0','1','0','1','0','1','0','0','1','0','0','0'),
            ('0','1','0','1','0','1','0','1','0','0','1','0','1','0'),
            ('0','1','0','1','0','1','0','1','0','0','1','1','0','0'),
            ('0','1','0','1','0','1','0','1','0','0','1','1','1','0'),
            ('0','1','0','1','0','1','0','1','0','1','0','0','0','0'),
            ('0','1','0','1','0','1','0','1','0','1','0','0','1','0'),
            ('0','1','0','1','0','1','0','1','0','1','0','1','0','0'),
            ('0','1','0','1','0','1','0','1','0','1','0','1','1','0'),
            ('0','1','0','1','0','1','0','1','0','1','1','0','0','0'),
            ('0','1','0','1','0','1','0','1','0','1','1','0','1','0'),
            ('0','1','0','1','0','1','0','1','0','1','1','1','0','0'),
            ('0','1','0','1','0','1','0','1','0','1','1','1','1','0'),
            ('0','1','0','1','0','1','0','1','1','0','0','0','0','0'),
            ('0','1','0','1','0','1','0','1','1','0','0','0','1','0'),
            ('0','1','0','1','0','1','0','1','1','0','0','1','0','0'),
            ('0','1','0','1','0','1','0','1','1','0','0','1','1','0'),
            ('0','1','0','1','0','1','0','1','1','0','1','0','0','0'),
            ('0','1','0','1','0','1','0','1','1','0','1','0','1','0'),
            ('0','1','0','1','0','1','0','1','1','0','1','1','0','0'),
            ('0','1','0','1','0','1','0','1','1','0','1','1','1','0'),
            ('0','1','0','1','0','1','0','1','1','1','0','0','0','0'),
            ('0','1','0','1','0','1','0','1','1','1','0','0','1','0'),
            ('0','1','0','1','0','1','0','1','1','1','0','1','0','0'),
            ('0','1','0','1','0','1','0','1','1','1','0','1','1','0'),
            ('0','1','0','1','0','1','0','1','1','1','1','0','0','0'),
            ('0','1','0','1','0','1','0','1','1','1','1','0','1','0'),
            ('0','1','0','1','0','1','0','1','1','1','1','1','0','0'),
            ('0','1','0','1','0','1','0','1','1','1','1','1','1','0'),
            ('0','1','0','1','0','1','1','0','0','0','0','0','0','0'),
            ('0','1','0','1','0','1','1','0','0','0','0','0','1','0'),
            ('0','1','0','1','0','1','1','0','0','0','0','1','0','0'),
            ('0','1','0','1','0','1','1','0','0','0','0','1','1','0'),
            ('0','1','0','1','0','1','1','0','0','0','1','0','0','0'),
            ('0','1','0','1','0','1','1','0','0','0','1','0','1','0'),
            ('0','1','0','1','0','1','1','0','0','0','1','1','0','0'),
            ('0','1','0','1','0','1','1','0','0','0','1','1','1','0'),
            ('0','1','0','1','0','1','1','0','0','1','0','0','0','0'),
            ('0','1','0','1','0','1','1','0','0','1','0','0','1','0'),
            ('0','1','0','1','0','1','1','0','0','1','0','1','0','0'),
            ('0','1','0','1','0','1','1','0','0','1','0','1','1','0'),
            ('0','1','0','1','0','1','1','0','0','1','1','0','0','0'),
            ('0','1','0','1','0','1','1','0','0','1','1','0','1','0'),
            ('0','1','0','1','0','1','1','0','0','1','1','1','0','0'),
            ('0','1','0','1','0','1','1','0','0','1','1','1','1','0'),
            ('0','1','0','1','0','1','1','0','1','0','0','0','0','0'),
            ('0','1','0','1','0','1','1','0','1','0','0','0','1','0'),
            ('0','1','0','1','0','1','1','0','1','0','0','1','0','0'),
            ('0','1','0','1','0','1','1','0','1','0','0','1','1','0'),
            ('0','1','0','1','0','1','1','0','1','0','1','0','0','0'),
            ('0','1','0','1','0','1','1','0','1','0','1','0','1','0'),
            ('0','1','0','1','0','1','1','0','1','0','1','1','0','0'),
            ('0','1','0','1','0','1','1','0','1','0','1','1','1','0'),
            ('0','1','0','1','0','1','1','0','1','1','0','0','0','0'),
            ('0','1','0','1','0','1','1','0','1','1','0','0','1','0'),
            ('0','1','0','1','0','1','1','0','1','1','0','1','0','0'),
            ('0','1','0','1','0','1','1','0','1','1','0','1','1','0'),
            ('0','1','0','1','0','1','1','0','1','1','1','0','0','0'),
            ('0','1','0','1','0','1','1','0','1','1','1','0','1','0'),
            ('0','1','0','1','0','1','1','0','1','1','1','1','0','0'),
            ('0','1','0','1','0','1','1','0','1','1','1','1','1','0'),
            ('0','1','0','1','0','1','1','1','0','0','0','0','0','0'),
            ('0','1','0','1','0','1','1','1','0','0','0','0','1','0'),
            ('0','1','0','1','0','1','1','1','0','0','0','1','0','0'),
            ('0','1','0','1','0','1','1','1','0','0','0','1','1','0'),
            ('0','1','0','1','0','1','1','1','0','0','1','0','0','0'),
            ('0','1','0','1','0','1','1','1','0','0','1','0','1','0'),
            ('0','1','0','1','0','1','1','1','0','0','1','1','0','0'),
            ('0','1','0','1','0','1','1','1','0','0','1','1','1','0'),
            ('0','1','0','1','0','1','1','1','0','1','0','0','0','0'),
            ('0','1','0','1','0','1','1','1','0','1','0','0','1','0'),
            ('0','1','0','1','0','1','1','1','0','1','0','1','0','0'),
            ('0','1','0','1','0','1','1','1','0','1','0','1','1','0'),
            ('0','1','0','1','0','1','1','1','0','1','1','0','0','0'),
            ('0','1','0','1','0','1','1','1','0','1','1','0','1','0'),
            ('0','1','0','1','0','1','1','1','0','1','1','1','0','0'),
            ('0','1','0','1','0','1','1','1','0','1','1','1','1','0'),
            ('0','1','0','1','0','1','1','1','1','0','0','0','0','0'),
            ('0','1','0','1','0','1','1','1','1','0','0','0','1','0'),
            ('0','1','0','1','0','1','1','1','1','0','0','1','0','0'),
            ('0','1','0','1','0','1','1','1','1','0','0','1','1','0'),
            ('0','1','0','1','0','1','1','1','1','0','1','0','0','0'),
            ('0','1','0','1','0','1','1','1','1','0','1','0','1','0'),
            ('0','1','0','1','0','1','1','1','1','0','1','1','0','0'),
            ('0','1','0','1','0','1','1','1','1','0','1','1','1','0'),
            ('0','1','0','1','0','1','1','1','1','1','0','0','0','0'),
            ('0','1','0','1','0','1','1','1','1','1','0','0','1','0'),
            ('0','1','0','1','0','1','1','1','1','1','0','1','0','0'),
            ('0','1','0','1','0','1','1','1','1','1','0','1','1','0'),
            ('0','1','0','1','0','1','1','1','1','1','1','0','0','0'),
            ('0','1','0','1','0','1','1','1','1','1','1','0','1','0'),
            ('0','1','0','1','0','1','1','1','1','1','1','1','0','0'),
            ('0','1','0','1','0','1','1','1','1','1','1','1','1','0'),
            ('0','1','0','1','1','0','0','0','0','0','0','0','0','0'),
            ('0','1','0','1','1','0','0','0','0','0','0','0','1','0'),
            ('0','1','0','1','1','0','0','0','0','0','0','1','0','0'),
            ('0','1','0','1','1','0','0','0','0','0','0','1','1','0'),
            ('0','1','0','1','1','0','0','0','0','0','1','0','0','0'),
            ('0','1','0','1','1','0','0','0','0','0','1','0','1','0'),
            ('0','1','0','1','1','0','0','0','0','0','1','1','0','0'),
            ('0','1','0','1','1','0','0','0','0','0','1','1','1','0'),
            ('0','1','0','1','1','0','0','0','0','1','0','0','0','0'),
            ('0','1','0','1','1','0','0','0','0','1','0','0','1','0'),
            ('0','1','0','1','1','0','0','0','0','1','0','1','0','0'),
            ('0','1','0','1','1','0','0','0','0','1','0','1','1','0'),
            ('0','1','0','1','1','0','0','0','0','1','1','0','0','0'),
            ('0','1','0','1','1','0','0','0','0','1','1','0','1','0'),
            ('0','1','0','1','1','0','0','0','0','1','1','1','0','0'),
            ('0','1','0','1','1','0','0','0','0','1','1','1','1','0'),
            ('0','1','0','1','1','0','0','0','1','0','0','0','0','0'),
            ('0','1','0','1','1','0','0','0','1','0','0','0','1','0'),
            ('0','1','0','1','1','0','0','0','1','0','0','1','0','0'),
            ('0','1','0','1','1','0','0','0','1','0','0','1','1','0'),
            ('0','1','0','1','1','0','0','0','1','0','1','0','0','0'),
            ('0','1','0','1','1','0','0','0','1','0','1','0','1','0'),
            ('0','1','0','1','1','0','0','0','1','0','1','1','0','0'),
            ('0','1','0','1','1','0','0','0','1','0','1','1','1','0'),
            ('0','1','0','1','1','0','0','0','1','1','0','0','0','0'),
            ('0','1','0','1','1','0','0','0','1','1','0','0','1','0'),
            ('0','1','0','1','1','0','0','0','1','1','0','1','0','0'),
            ('0','1','0','1','1','0','0','0','1','1','0','1','1','0'),
            ('0','1','0','1','1','0','0','0','1','1','1','0','0','0'),
            ('0','1','0','1','1','0','0','0','1','1','1','0','1','0'),
            ('0','1','0','1','1','0','0','0','1','1','1','1','0','0'),
            ('0','1','0','1','1','0','0','0','1','1','1','1','1','0'),
            ('0','1','0','1','1','0','0','1','0','0','0','0','0','0'),
            ('0','1','0','1','1','0','0','1','0','0','0','0','1','0'),
            ('0','1','0','1','1','0','0','1','0','0','0','1','0','0'),
            ('0','1','0','1','1','0','0','1','0','0','0','1','1','0'),
            ('0','1','0','1','1','0','0','1','0','0','1','0','0','0'),
            ('0','1','0','1','1','0','0','1','0','0','1','0','1','0'),
            ('0','1','0','1','1','0','0','1','0','0','1','1','0','0'),
            ('0','1','0','1','1','0','0','1','0','0','1','1','1','0'),
            ('0','1','0','1','1','0','0','1','0','1','0','0','0','0'),
            ('0','1','0','1','1','0','0','1','0','1','0','0','1','0'),
            ('0','1','0','1','1','0','0','1','0','1','0','1','0','0'),
            ('0','1','0','1','1','0','0','1','0','1','0','1','1','0'),
            ('0','1','0','1','1','0','0','1','0','1','1','0','0','0'),
            ('0','1','0','1','1','0','0','1','0','1','1','0','1','0'),
            ('0','1','0','1','1','0','0','1','0','1','1','1','0','0'),
            ('0','1','0','1','1','0','0','1','0','1','1','1','1','0'),
            ('0','1','0','1','1','0','0','1','1','0','0','0','0','0'),
            ('0','1','0','1','1','0','0','1','1','0','0','0','1','0'),
            ('0','1','0','1','1','0','0','1','1','0','0','1','0','0'),
            ('0','1','0','1','1','0','0','1','1','0','0','1','1','0'),
            ('0','1','0','1','1','0','0','1','1','0','1','0','0','0'),
            ('0','1','0','1','1','0','0','1','1','0','1','0','1','0'),
            ('0','1','0','1','1','0','0','1','1','0','1','1','0','0'),
            ('0','1','0','1','1','0','0','1','1','0','1','1','1','0'),
            ('0','1','0','1','1','0','0','1','1','1','0','0','0','0'),
            ('0','1','0','1','1','0','0','1','1','1','0','0','1','0'),
            ('0','1','0','1','1','0','0','1','1','1','0','1','0','0'),
            ('0','1','0','1','1','0','0','1','1','1','0','1','1','0'),
            ('0','1','0','1','1','0','0','1','1','1','1','0','0','0'),
            ('0','1','0','1','1','0','0','1','1','1','1','0','1','0'),
            ('0','1','0','1','1','0','0','1','1','1','1','1','0','0'),
            ('0','1','0','1','1','0','0','1','1','1','1','1','1','0'),
            ('0','1','0','1','1','0','1','0','0','0','0','0','0','0'),
            ('0','1','0','1','1','0','1','0','0','0','0','0','1','0'),
            ('0','1','0','1','1','0','1','0','0','0','0','1','0','0'),
            ('0','1','0','1','1','0','1','0','0','0','0','1','1','0'),
            ('0','1','0','1','1','0','1','0','0','0','1','0','0','0'),
            ('0','1','0','1','1','0','1','0','0','0','1','0','1','0'),
            ('0','1','0','1','1','0','1','0','0','0','1','1','0','0'),
            ('0','1','0','1','1','0','1','0','0','0','1','1','1','0'),
            ('0','1','0','1','1','0','1','0','0','1','0','0','0','0'),
            ('0','1','0','1','1','0','1','0','0','1','0','0','1','0'),
            ('0','1','0','1','1','0','1','0','0','1','0','1','0','0'),
            ('0','1','0','1','1','0','1','0','0','1','0','1','1','0'),
            ('0','1','0','1','1','0','1','0','0','1','1','0','0','0'),
            ('0','1','0','1','1','0','1','0','0','1','1','0','1','0'),
            ('0','1','0','1','1','0','1','0','0','1','1','1','0','0'),
            ('0','1','0','1','1','0','1','0','0','1','1','1','1','0'),
            ('0','1','0','1','1','0','1','0','1','0','0','0','0','0'),
            ('0','1','0','1','1','0','1','0','1','0','0','0','1','0'),
            ('0','1','0','1','1','0','1','0','1','0','0','1','0','0'),
            ('0','1','0','1','1','0','1','0','1','0','0','1','1','0'),
            ('0','1','0','1','1','0','1','0','1','0','1','0','0','0'),
            ('0','1','0','1','1','0','1','0','1','0','1','0','1','0'),
            ('0','1','0','1','1','0','1','0','1','0','1','1','0','0'),
            ('0','1','0','1','1','0','1','0','1','0','1','1','1','0'),
            ('0','1','0','1','1','0','1','0','1','1','0','0','0','0'),
            ('0','1','0','1','1','0','1','0','1','1','0','0','1','0'),
            ('0','1','0','1','1','0','1','0','1','1','0','1','0','0'),
            ('0','1','0','1','1','0','1','0','1','1','0','1','1','0'),
            ('0','1','0','1','1','0','1','0','1','1','1','0','0','0'),
            ('0','1','0','1','1','0','1','0','1','1','1','0','1','0'),
            ('0','1','0','1','1','0','1','0','1','1','1','1','0','0'),
            ('0','1','0','1','1','0','1','0','1','1','1','1','1','0'),
            ('0','1','0','1','1','0','1','1','0','0','0','0','0','0'),
            ('0','1','0','1','1','0','1','1','0','0','0','0','1','0'),
            ('0','1','0','1','1','0','1','1','0','0','0','1','0','0'),
            ('0','1','0','1','1','0','1','1','0','0','0','1','1','0'),
            ('0','1','0','1','1','0','1','1','0','0','1','0','0','0'),
            ('0','1','0','1','1','0','1','1','0','0','1','0','1','0'),
            ('0','1','0','1','1','0','1','1','0','0','1','1','0','0'),
            ('0','1','0','1','1','0','1','1','0','0','1','1','1','0'),
            ('0','1','0','1','1','0','1','1','0','1','0','0','0','0'),
            ('0','1','0','1','1','0','1','1','0','1','0','0','1','0'),
            ('0','1','0','1','1','0','1','1','0','1','0','1','0','0'),
            ('0','1','0','1','1','0','1','1','0','1','0','1','1','0'),
            ('0','1','0','1','1','0','1','1','0','1','1','0','0','0'),
            ('0','1','0','1','1','0','1','1','0','1','1','0','1','0'),
            ('0','1','0','1','1','0','1','1','0','1','1','1','0','0'),
            ('0','1','0','1','1','0','1','1','0','1','1','1','1','0'),
            ('0','1','0','1','1','0','1','1','1','0','0','0','0','0'),
            ('0','1','0','1','1','0','1','1','1','0','0','0','1','0'),
            ('0','1','0','1','1','0','1','1','1','0','0','1','0','0'),
            ('0','1','0','1','1','0','1','1','1','0','0','1','1','0'),
            ('0','1','0','1','1','0','1','1','1','0','1','0','0','0'),
            ('0','1','0','1','1','0','1','1','1','0','1','0','1','0'),
            ('0','1','0','1','1','0','1','1','1','0','1','1','0','0'),
            ('0','1','0','1','1','0','1','1','1','0','1','1','1','0'),
            ('0','1','0','1','1','0','1','1','1','1','0','0','0','0'),
            ('0','1','0','1','1','0','1','1','1','1','0','0','1','0'),
            ('0','1','0','1','1','0','1','1','1','1','0','1','0','0'),
            ('0','1','0','1','1','0','1','1','1','1','0','1','1','0'),
            ('0','1','0','1','1','0','1','1','1','1','1','0','0','0'),
            ('0','1','0','1','1','0','1','1','1','1','1','0','1','0'),
            ('0','1','0','1','1','0','1','1','1','1','1','1','0','0'),
            ('0','1','0','1','1','0','1','1','1','1','1','1','1','0'),
            ('0','1','0','1','1','1','0','0','0','0','0','0','0','0'),
            ('0','1','0','1','1','1','0','0','0','0','0','0','1','0'),
            ('0','1','0','1','1','1','0','0','0','0','0','1','0','0'),
            ('0','1','0','1','1','1','0','0','0','0','0','1','1','0'),
            ('0','1','0','1','1','1','0','0','0','0','1','0','0','0'),
            ('0','1','0','1','1','1','0','0','0','0','1','0','1','0'),
            ('0','1','0','1','1','1','0','0','0','0','1','1','0','0'),
            ('0','1','0','1','1','1','0','0','0','0','1','1','1','0'),
            ('0','1','0','1','1','1','0','0','0','1','0','0','0','0'),
            ('0','1','0','1','1','1','0','0','0','1','0','0','1','0'),
            ('0','1','0','1','1','1','0','0','0','1','0','1','0','0'),
            ('0','1','0','1','1','1','0','0','0','1','0','1','1','0'),
            ('0','1','0','1','1','1','0','0','0','1','1','0','0','0'),
            ('0','1','0','1','1','1','0','0','0','1','1','0','1','0'),
            ('0','1','0','1','1','1','0','0','0','1','1','1','0','0'),
            ('0','1','0','1','1','1','0','0','0','1','1','1','1','0'),
            ('0','1','0','1','1','1','0','0','1','0','0','0','0','0'),
            ('0','1','0','1','1','1','0','0','1','0','0','0','1','0'),
            ('0','1','0','1','1','1','0','0','1','0','0','1','0','0'),
            ('0','1','0','1','1','1','0','0','1','0','0','1','1','0'),
            ('0','1','0','1','1','1','0','0','1','0','1','0','0','0'),
            ('0','1','0','1','1','1','0','0','1','0','1','0','1','0'),
            ('0','1','0','1','1','1','0','0','1','0','1','1','0','0'),
            ('0','1','0','1','1','1','0','0','1','0','1','1','1','0'),
            ('0','1','0','1','1','1','0','0','1','1','0','0','0','0'),
            ('0','1','0','1','1','1','0','0','1','1','0','0','1','0'),
            ('0','1','0','1','1','1','0','0','1','1','0','1','0','0'),
            ('0','1','0','1','1','1','0','0','1','1','0','1','1','0'),
            ('0','1','0','1','1','1','0','0','1','1','1','0','0','0'),
            ('0','1','0','1','1','1','0','0','1','1','1','0','1','0'),
            ('0','1','0','1','1','1','0','0','1','1','1','1','0','0'),
            ('0','1','0','1','1','1','0','0','1','1','1','1','1','0'),
            ('0','1','0','1','1','1','0','1','0','0','0','0','0','0'),
            ('0','1','0','1','1','1','0','1','0','0','0','0','1','0'),
            ('0','1','0','1','1','1','0','1','0','0','0','1','0','0'),
            ('0','1','0','1','1','1','0','1','0','0','0','1','1','0'),
            ('0','1','0','1','1','1','0','1','0','0','1','0','0','0'),
            ('0','1','0','1','1','1','0','1','0','0','1','0','1','0'),
            ('0','1','0','1','1','1','0','1','0','0','1','1','0','0'),
            ('0','1','0','1','1','1','0','1','0','0','1','1','1','0'),
            ('0','1','0','1','1','1','0','1','0','1','0','0','0','0'),
            ('0','1','0','1','1','1','0','1','0','1','0','0','1','0'),
            ('0','1','0','1','1','1','0','1','0','1','0','1','0','0'),
            ('0','1','0','1','1','1','0','1','0','1','0','1','1','0'),
            ('0','1','0','1','1','1','0','1','0','1','1','0','0','0'),
            ('0','1','0','1','1','1','0','1','0','1','1','0','1','0'),
            ('0','1','0','1','1','1','0','1','0','1','1','1','0','0'),
            ('0','1','0','1','1','1','0','1','0','1','1','1','1','0'),
            ('0','1','0','1','1','1','0','1','1','0','0','0','0','0'),
            ('0','1','0','1','1','1','0','1','1','0','0','0','1','0'),
            ('0','1','0','1','1','1','0','1','1','0','0','1','0','0'),
            ('0','1','0','1','1','1','0','1','1','0','0','1','1','0'),
            ('0','1','0','1','1','1','0','1','1','0','1','0','0','0'),
            ('0','1','0','1','1','1','0','1','1','0','1','0','1','0'),
            ('0','1','0','1','1','1','0','1','1','0','1','1','0','0'),
            ('0','1','0','1','1','1','0','1','1','0','1','1','1','0'),
            ('0','1','0','1','1','1','0','1','1','1','0','0','0','0'),
            ('0','1','0','1','1','1','0','1','1','1','0','0','1','0'),
            ('0','1','0','1','1','1','0','1','1','1','0','1','0','0'),
            ('0','1','0','1','1','1','0','1','1','1','0','1','1','0'),
            ('0','1','0','1','1','1','0','1','1','1','1','0','0','0'),
            ('0','1','0','1','1','1','0','1','1','1','1','0','1','0'),
            ('0','1','0','1','1','1','0','1','1','1','1','1','0','0'),
            ('0','1','0','1','1','1','0','1','1','1','1','1','1','0'),
            ('0','1','0','1','1','1','1','0','0','0','0','0','0','0'),
            ('0','1','0','1','1','1','1','0','0','0','0','0','1','0'),
            ('0','1','0','1','1','1','1','0','0','0','0','1','0','0'),
            ('0','1','0','1','1','1','1','0','0','0','0','1','1','0'),
            ('0','1','0','1','1','1','1','0','0','0','1','0','0','0'),
            ('0','1','0','1','1','1','1','0','0','0','1','0','1','0'),
            ('0','1','0','1','1','1','1','0','0','0','1','1','0','0'),
            ('0','1','0','1','1','1','1','0','0','0','1','1','1','0'),
            ('0','1','0','1','1','1','1','0','0','1','0','0','0','0'),
            ('0','1','0','1','1','1','1','0','0','1','0','0','1','0'),
            ('0','1','0','1','1','1','1','0','0','1','0','1','0','0'),
            ('0','1','0','1','1','1','1','0','0','1','0','1','1','0'),
            ('0','1','0','1','1','1','1','0','0','1','1','0','0','0'),
            ('0','1','0','1','1','1','1','0','0','1','1','0','1','0'),
            ('0','1','0','1','1','1','1','0','0','1','1','1','0','0'),
            ('0','1','0','1','1','1','1','0','0','1','1','1','1','0'),
            ('0','1','0','1','1','1','1','0','1','0','0','0','0','0'),
            ('0','1','0','1','1','1','1','0','1','0','0','0','1','0'),
            ('0','1','0','1','1','1','1','0','1','0','0','1','0','0'),
            ('0','1','0','1','1','1','1','0','1','0','0','1','1','0'),
            ('0','1','0','1','1','1','1','0','1','0','1','0','0','0'),
            ('0','1','0','1','1','1','1','0','1','0','1','0','1','0'),
            ('0','1','0','1','1','1','1','0','1','0','1','1','0','0'),
            ('0','1','0','1','1','1','1','0','1','0','1','1','1','0'),
            ('0','1','0','1','1','1','1','0','1','1','0','0','0','0'),
            ('0','1','0','1','1','1','1','0','1','1','0','0','1','0'),
            ('0','1','0','1','1','1','1','0','1','1','0','1','0','0'),
            ('0','1','0','1','1','1','1','0','1','1','0','1','1','0'),
            ('0','1','0','1','1','1','1','0','1','1','1','0','0','0'),
            ('0','1','0','1','1','1','1','0','1','1','1','0','1','0'),
            ('0','1','0','1','1','1','1','0','1','1','1','1','0','0'),
            ('0','1','0','1','1','1','1','0','1','1','1','1','1','0'),
            ('0','1','0','1','1','1','1','1','0','0','0','0','0','0'),
            ('0','1','0','1','1','1','1','1','0','0','0','0','1','0'),
            ('0','1','0','1','1','1','1','1','0','0','0','1','0','0'),
            ('0','1','0','1','1','1','1','1','0','0','0','1','1','0'),
            ('0','1','0','1','1','1','1','1','0','0','1','0','0','0'),
            ('0','1','0','1','1','1','1','1','0','0','1','0','1','0'),
            ('0','1','0','1','1','1','1','1','0','0','1','1','0','0'),
            ('0','1','0','1','1','1','1','1','0','0','1','1','1','0'),
            ('0','1','0','1','1','1','1','1','0','1','0','0','0','0'),
            ('0','1','0','1','1','1','1','1','0','1','0','0','1','0'),
            ('0','1','0','1','1','1','1','1','0','1','0','1','0','0'),
            ('0','1','0','1','1','1','1','1','0','1','0','1','1','0'),
            ('0','1','0','1','1','1','1','1','0','1','1','0','0','0'),
            ('0','1','0','1','1','1','1','1','0','1','1','0','1','0'),
            ('0','1','0','1','1','1','1','1','0','1','1','1','0','0'),
            ('0','1','0','1','1','1','1','1','0','1','1','1','1','0'),
            ('0','1','0','1','1','1','1','1','1','0','0','0','0','0'),
            ('0','1','0','1','1','1','1','1','1','0','0','0','1','0'),
            ('0','1','0','1','1','1','1','1','1','0','0','1','0','0'),
            ('0','1','0','1','1','1','1','1','1','0','0','1','1','0'),
            ('0','1','0','1','1','1','1','1','1','0','1','0','0','0'),
            ('0','1','0','1','1','1','1','1','1','0','1','0','1','0'),
            ('0','1','0','1','1','1','1','1','1','0','1','1','0','0'),
            ('0','1','0','1','1','1','1','1','1','0','1','1','1','0'),
            ('0','1','0','1','1','1','1','1','1','1','0','0','0','0'),
            ('0','1','0','1','1','1','1','1','1','1','0','0','1','0'),
            ('0','1','0','1','1','1','1','1','1','1','0','1','0','0'),
            ('0','1','0','1','1','1','1','1','1','1','0','1','1','0'),
            ('0','1','0','1','1','1','1','1','1','1','1','0','0','0'),
            ('0','1','0','1','1','1','1','1','1','1','1','0','1','0'),
            ('0','1','0','1','1','1','1','1','1','1','1','1','0','0'),
            ('0','1','0','1','1','1','1','1','1','1','1','1','1','0'),
            ('0','1','1','0','0','0','0','0','0','0','0','0','0','0'),
            ('0','1','1','0','0','0','0','0','0','0','0','0','1','0'),
            ('0','1','1','0','0','0','0','0','0','0','0','1','0','0'),
            ('0','1','1','0','0','0','0','0','0','0','0','1','1','0'),
            ('0','1','1','0','0','0','0','0','0','0','1','0','0','0'),
            ('0','1','1','0','0','0','0','0','0','0','1','0','1','0'),
            ('0','1','1','0','0','0','0','0','0','0','1','1','0','0'),
            ('0','1','1','0','0','0','0','0','0','0','1','1','1','0'),
            ('0','1','1','0','0','0','0','0','0','1','0','0','0','0'),
            ('0','1','1','0','0','0','0','0','0','1','0','0','1','0'),
            ('0','1','1','0','0','0','0','0','0','1','0','1','0','0'),
            ('0','1','1','0','0','0','0','0','0','1','0','1','1','0'),
            ('0','1','1','0','0','0','0','0','0','1','1','0','0','0'),
            ('0','1','1','0','0','0','0','0','0','1','1','0','1','0'),
            ('0','1','1','0','0','0','0','0','0','1','1','1','0','0'),
            ('0','1','1','0','0','0','0','0','0','1','1','1','1','0'),
            ('0','1','1','0','0','0','0','0','1','0','0','0','0','0'),
            ('0','1','1','0','0','0','0','0','1','0','0','0','1','0'),
            ('0','1','1','0','0','0','0','0','1','0','0','1','0','0'),
            ('0','1','1','0','0','0','0','0','1','0','0','1','1','0'),
            ('0','1','1','0','0','0','0','0','1','0','1','0','0','0'),
            ('0','1','1','0','0','0','0','0','1','0','1','0','1','0'),
            ('0','1','1','0','0','0','0','0','1','0','1','1','0','0'),
            ('0','1','1','0','0','0','0','0','1','0','1','1','1','0'),
            ('0','1','1','0','0','0','0','0','1','1','0','0','0','0'),
            ('0','1','1','0','0','0','0','0','1','1','0','0','1','0'),
            ('0','1','1','0','0','0','0','0','1','1','0','1','0','0'),
            ('0','1','1','0','0','0','0','0','1','1','0','1','1','0'),
            ('0','1','1','0','0','0','0','0','1','1','1','0','0','0'),
            ('0','1','1','0','0','0','0','0','1','1','1','0','1','0'),
            ('0','1','1','0','0','0','0','0','1','1','1','1','0','0'),
            ('0','1','1','0','0','0','0','0','1','1','1','1','1','0'),
            ('0','1','1','0','0','0','0','1','0','0','0','0','0','0'),
            ('0','1','1','0','0','0','0','1','0','0','0','0','1','0'),
            ('0','1','1','0','0','0','0','1','0','0','0','1','0','0'),
            ('0','1','1','0','0','0','0','1','0','0','0','1','1','0'),
            ('0','1','1','0','0','0','0','1','0','0','1','0','0','0'),
            ('0','1','1','0','0','0','0','1','0','0','1','0','1','0'),
            ('0','1','1','0','0','0','0','1','0','0','1','1','0','0'),
            ('0','1','1','0','0','0','0','1','0','0','1','1','1','0'),
            ('0','1','1','0','0','0','0','1','0','1','0','0','0','0'),
            ('0','1','1','0','0','0','0','1','0','1','0','0','1','0'),
            ('0','1','1','0','0','0','0','1','0','1','0','1','0','0'),
            ('0','1','1','0','0','0','0','1','0','1','0','1','1','0'),
            ('0','1','1','0','0','0','0','1','0','1','1','0','0','0'),
            ('0','1','1','0','0','0','0','1','0','1','1','0','1','0'),
            ('0','1','1','0','0','0','0','1','0','1','1','1','0','0'),
            ('0','1','1','0','0','0','0','1','0','1','1','1','1','0'),
            ('0','1','1','0','0','0','0','1','1','0','0','0','0','0'),
            ('0','1','1','0','0','0','0','1','1','0','0','0','1','0'),
            ('0','1','1','0','0','0','0','1','1','0','0','1','0','0'),
            ('0','1','1','0','0','0','0','1','1','0','0','1','1','0'),
            ('0','1','1','0','0','0','0','1','1','0','1','0','0','0'),
            ('0','1','1','0','0','0','0','1','1','0','1','0','1','0'),
            ('0','1','1','0','0','0','0','1','1','0','1','1','0','0'),
            ('0','1','1','0','0','0','0','1','1','0','1','1','1','0'),
            ('0','1','1','0','0','0','0','1','1','1','0','0','0','0'),
            ('0','1','1','0','0','0','0','1','1','1','0','0','1','0'),
            ('0','1','1','0','0','0','0','1','1','1','0','1','0','0'),
            ('0','1','1','0','0','0','0','1','1','1','0','1','1','0'),
            ('0','1','1','0','0','0','0','1','1','1','1','0','0','0'),
            ('0','1','1','0','0','0','0','1','1','1','1','0','1','0'),
            ('0','1','1','0','0','0','0','1','1','1','1','1','0','0'),
            ('0','1','1','0','0','0','0','1','1','1','1','1','1','0'),
            ('0','1','1','0','0','0','1','0','0','0','0','0','0','0'),
            ('0','1','1','0','0','0','1','0','0','0','0','0','1','0'),
            ('0','1','1','0','0','0','1','0','0','0','0','1','0','0'),
            ('0','1','1','0','0','0','1','0','0','0','0','1','1','0'),
            ('0','1','1','0','0','0','1','0','0','0','1','0','0','0'),
            ('0','1','1','0','0','0','1','0','0','0','1','0','1','0'),
            ('0','1','1','0','0','0','1','0','0','0','1','1','0','0'),
            ('0','1','1','0','0','0','1','0','0','0','1','1','1','0'),
            ('0','1','1','0','0','0','1','0','0','1','0','0','0','0'),
            ('0','1','1','0','0','0','1','0','0','1','0','0','1','0'),
            ('0','1','1','0','0','0','1','0','0','1','0','1','0','0'),
            ('0','1','1','0','0','0','1','0','0','1','0','1','1','0'),
            ('0','1','1','0','0','0','1','0','0','1','1','0','0','0'),
            ('0','1','1','0','0','0','1','0','0','1','1','0','1','0'),
            ('0','1','1','0','0','0','1','0','0','1','1','1','0','0'),
            ('0','1','1','0','0','0','1','0','0','1','1','1','1','0'),
            ('0','1','1','0','0','0','1','0','1','0','0','0','0','0'),
            ('0','1','1','0','0','0','1','0','1','0','0','0','1','0'),
            ('0','1','1','0','0','0','1','0','1','0','0','1','0','0'),
            ('0','1','1','0','0','0','1','0','1','0','0','1','1','0'),
            ('0','1','1','0','0','0','1','0','1','0','1','0','0','0'),
            ('0','1','1','0','0','0','1','0','1','0','1','0','1','0'),
            ('0','1','1','0','0','0','1','0','1','0','1','1','0','0'),
            ('0','1','1','0','0','0','1','0','1','0','1','1','1','0'),
            ('0','1','1','0','0','0','1','0','1','1','0','0','0','0'),
            ('0','1','1','0','0','0','1','0','1','1','0','0','1','0'),
            ('0','1','1','0','0','0','1','0','1','1','0','1','0','0'),
            ('0','1','1','0','0','0','1','0','1','1','0','1','1','0'),
            ('0','1','1','0','0','0','1','0','1','1','1','0','0','0'),
            ('0','1','1','0','0','0','1','0','1','1','1','0','1','0'),
            ('0','1','1','0','0','0','1','0','1','1','1','1','0','0'),
            ('0','1','1','0','0','0','1','0','1','1','1','1','1','0'),
            ('0','1','1','0','0','0','1','1','0','0','0','0','0','0'),
            ('0','1','1','0','0','0','1','1','0','0','0','0','1','0'),
            ('0','1','1','0','0','0','1','1','0','0','0','1','0','0'),
            ('0','1','1','0','0','0','1','1','0','0','0','1','1','0'),
            ('0','1','1','0','0','0','1','1','0','0','1','0','0','0'),
            ('0','1','1','0','0','0','1','1','0','0','1','0','1','0'),
            ('0','1','1','0','0','0','1','1','0','0','1','1','0','0'),
            ('0','1','1','0','0','0','1','1','0','0','1','1','1','0'),
            ('0','1','1','0','0','0','1','1','0','1','0','0','0','0'),
            ('0','1','1','0','0','0','1','1','0','1','0','0','1','0'),
            ('0','1','1','0','0','0','1','1','0','1','0','1','0','0'),
            ('0','1','1','0','0','0','1','1','0','1','0','1','1','0'),
            ('0','1','1','0','0','0','1','1','0','1','1','0','0','0'),
            ('0','1','1','0','0','0','1','1','0','1','1','0','1','0'),
            ('0','1','1','0','0','0','1','1','0','1','1','1','0','0'),
            ('0','1','1','0','0','0','1','1','0','1','1','1','1','0'),
            ('0','1','1','0','0','0','1','1','1','0','0','0','0','0'),
            ('0','1','1','0','0','0','1','1','1','0','0','0','1','0'),
            ('0','1','1','0','0','0','1','1','1','0','0','1','0','0'),
            ('0','1','1','0','0','0','1','1','1','0','0','1','1','0'),
            ('0','1','1','0','0','0','1','1','1','0','1','0','0','0'),
            ('0','1','1','0','0','0','1','1','1','0','1','0','1','0'),
            ('0','1','1','0','0','0','1','1','1','0','1','1','0','0'),
            ('0','1','1','0','0','0','1','1','1','0','1','1','1','0'),
            ('0','1','1','0','0','0','1','1','1','1','0','0','0','0'),
            ('0','1','1','0','0','0','1','1','1','1','0','0','1','0'),
            ('0','1','1','0','0','0','1','1','1','1','0','1','0','0'),
            ('0','1','1','0','0','0','1','1','1','1','0','1','1','0'),
            ('0','1','1','0','0','0','1','1','1','1','1','0','0','0'),
            ('0','1','1','0','0','0','1','1','1','1','1','0','1','0'),
            ('0','1','1','0','0','0','1','1','1','1','1','1','0','0'),
            ('0','1','1','0','0','0','1','1','1','1','1','1','1','0'),
            ('0','1','1','0','0','1','0','0','0','0','0','0','0','0'),
            ('0','1','1','0','0','1','0','0','0','0','0','0','1','0'),
            ('0','1','1','0','0','1','0','0','0','0','0','1','0','0'),
            ('0','1','1','0','0','1','0','0','0','0','0','1','1','0'),
            ('0','1','1','0','0','1','0','0','0','0','1','0','0','0'),
            ('0','1','1','0','0','1','0','0','0','0','1','0','1','0'),
            ('0','1','1','0','0','1','0','0','0','0','1','1','0','0'),
            ('0','1','1','0','0','1','0','0','0','0','1','1','1','0'),
            ('0','1','1','0','0','1','0','0','0','1','0','0','0','0'),
            ('0','1','1','0','0','1','0','0','0','1','0','0','1','0'),
            ('0','1','1','0','0','1','0','0','0','1','0','1','0','0'),
            ('0','1','1','0','0','1','0','0','0','1','0','1','1','0'),
            ('0','1','1','0','0','1','0','0','0','1','1','0','0','0'),
            ('0','1','1','0','0','1','0','0','0','1','1','0','1','0'),
            ('0','1','1','0','0','1','0','0','0','1','1','1','0','0'),
            ('0','1','1','0','0','1','0','0','0','1','1','1','1','0'),
            ('0','1','1','0','0','1','0','0','1','0','0','0','0','0'),
            ('0','1','1','0','0','1','0','0','1','0','0','0','1','0'),
            ('0','1','1','0','0','1','0','0','1','0','0','1','0','0'),
            ('0','1','1','0','0','1','0','0','1','0','0','1','1','0'),
            ('0','1','1','0','0','1','0','0','1','0','1','0','0','0'),
            ('0','1','1','0','0','1','0','0','1','0','1','0','1','0'),
            ('0','1','1','0','0','1','0','0','1','0','1','1','0','0'),
            ('0','1','1','0','0','1','0','0','1','0','1','1','1','0'),
            ('0','1','1','0','0','1','0','0','1','1','0','0','0','0'),
            ('0','1','1','0','0','1','0','0','1','1','0','0','1','0'),
            ('0','1','1','0','0','1','0','0','1','1','0','1','0','0'),
            ('0','1','1','0','0','1','0','0','1','1','0','1','1','0'),
            ('0','1','1','0','0','1','0','0','1','1','1','0','0','0'),
            ('0','1','1','0','0','1','0','0','1','1','1','0','1','0'),
            ('0','1','1','0','0','1','0','0','1','1','1','1','0','0'),
            ('0','1','1','0','0','1','0','0','1','1','1','1','1','0'),
            ('0','1','1','0','0','1','0','1','0','0','0','0','0','0'),
            ('0','1','1','0','0','1','0','1','0','0','0','0','1','0'),
            ('0','1','1','0','0','1','0','1','0','0','0','1','0','0'),
            ('0','1','1','0','0','1','0','1','0','0','0','1','1','0'),
            ('0','1','1','0','0','1','0','1','0','0','1','0','0','0'),
            ('0','1','1','0','0','1','0','1','0','0','1','0','1','0'),
            ('0','1','1','0','0','1','0','1','0','0','1','1','0','0'),
            ('0','1','1','0','0','1','0','1','0','0','1','1','1','0'),
            ('0','1','1','0','0','1','0','1','0','1','0','0','0','0'),
            ('0','1','1','0','0','1','0','1','0','1','0','0','1','0'),
            ('0','1','1','0','0','1','0','1','0','1','0','1','0','0'),
            ('0','1','1','0','0','1','0','1','0','1','0','1','1','0'),
            ('0','1','1','0','0','1','0','1','0','1','1','0','0','0'),
            ('0','1','1','0','0','1','0','1','0','1','1','0','1','0'),
            ('0','1','1','0','0','1','0','1','0','1','1','1','0','0'),
            ('0','1','1','0','0','1','0','1','0','1','1','1','1','0'),
            ('0','1','1','0','0','1','0','1','1','0','0','0','0','0'),
            ('0','1','1','0','0','1','0','1','1','0','0','0','1','0'),
            ('0','1','1','0','0','1','0','1','1','0','0','1','0','0'),
            ('0','1','1','0','0','1','0','1','1','0','0','1','1','0'),
            ('0','1','1','0','0','1','0','1','1','0','1','0','0','0'),
            ('0','1','1','0','0','1','0','1','1','0','1','0','1','0'),
            ('0','1','1','0','0','1','0','1','1','0','1','1','0','0'),
            ('0','1','1','0','0','1','0','1','1','0','1','1','1','0'),
            ('0','1','1','0','0','1','0','1','1','1','0','0','0','0'),
            ('0','1','1','0','0','1','0','1','1','1','0','0','1','0'),
            ('0','1','1','0','0','1','0','1','1','1','0','1','0','0'),
            ('0','1','1','0','0','1','0','1','1','1','0','1','1','0'),
            ('0','1','1','0','0','1','0','1','1','1','1','0','0','0'),
            ('0','1','1','0','0','1','0','1','1','1','1','0','1','0'),
            ('0','1','1','0','0','1','0','1','1','1','1','1','0','0'),
            ('0','1','1','0','0','1','0','1','1','1','1','1','1','0'),
            ('0','1','1','0','0','1','1','0','0','0','0','0','0','0'),
            ('0','1','1','0','0','1','1','0','0','0','0','0','1','0'),
            ('0','1','1','0','0','1','1','0','0','0','0','1','0','0'),
            ('0','1','1','0','0','1','1','0','0','0','0','1','1','0'),
            ('0','1','1','0','0','1','1','0','0','0','1','0','0','0'),
            ('0','1','1','0','0','1','1','0','0','0','1','0','1','0'),
            ('0','1','1','0','0','1','1','0','0','0','1','1','0','0'),
            ('0','1','1','0','0','1','1','0','0','0','1','1','1','0'),
            ('0','1','1','0','0','1','1','0','0','1','0','0','0','0'),
            ('0','1','1','0','0','1','1','0','0','1','0','0','1','0'),
            ('0','1','1','0','0','1','1','0','0','1','0','1','0','0'),
            ('0','1','1','0','0','1','1','0','0','1','0','1','1','0'),
            ('0','1','1','0','0','1','1','0','0','1','1','0','0','0'),
            ('0','1','1','0','0','1','1','0','0','1','1','0','1','0'),
            ('0','1','1','0','0','1','1','0','0','1','1','1','0','0'),
            ('0','1','1','0','0','1','1','0','0','1','1','1','1','0'),
            ('0','1','1','0','0','1','1','0','1','0','0','0','0','0'),
            ('0','1','1','0','0','1','1','0','1','0','0','0','1','0'),
            ('0','1','1','0','0','1','1','0','1','0','0','1','0','0'),
            ('0','1','1','0','0','1','1','0','1','0','0','1','1','0'),
            ('0','1','1','0','0','1','1','0','1','0','1','0','0','0'),
            ('0','1','1','0','0','1','1','0','1','0','1','0','1','0'),
            ('0','1','1','0','0','1','1','0','1','0','1','1','0','0'),
            ('0','1','1','0','0','1','1','0','1','0','1','1','1','0'),
            ('0','1','1','0','0','1','1','0','1','1','0','0','0','0'),
            ('0','1','1','0','0','1','1','0','1','1','0','0','1','0'),
            ('0','1','1','0','0','1','1','0','1','1','0','1','0','0'),
            ('0','1','1','0','0','1','1','0','1','1','0','1','1','0'),
            ('0','1','1','0','0','1','1','0','1','1','1','0','0','0'),
            ('0','1','1','0','0','1','1','0','1','1','1','0','1','0'),
            ('0','1','1','0','0','1','1','0','1','1','1','1','0','0'),
            ('0','1','1','0','0','1','1','0','1','1','1','1','1','0'),
            ('0','1','1','0','0','1','1','1','0','0','0','0','0','0'),
            ('0','1','1','0','0','1','1','1','0','0','0','0','1','0'),
            ('0','1','1','0','0','1','1','1','0','0','0','1','0','0'),
            ('0','1','1','0','0','1','1','1','0','0','0','1','1','0'),
            ('0','1','1','0','0','1','1','1','0','0','1','0','0','0'),
            ('0','1','1','0','0','1','1','1','0','0','1','0','1','0'),
            ('0','1','1','0','0','1','1','1','0','0','1','1','0','0'),
            ('0','1','1','0','0','1','1','1','0','0','1','1','1','0'),
            ('0','1','1','0','0','1','1','1','0','1','0','0','0','0'),
            ('0','1','1','0','0','1','1','1','0','1','0','0','1','0'),
            ('0','1','1','0','0','1','1','1','0','1','0','1','0','0'),
            ('0','1','1','0','0','1','1','1','0','1','0','1','1','0'),
            ('0','1','1','0','0','1','1','1','0','1','1','0','0','0'),
            ('0','1','1','0','0','1','1','1','0','1','1','0','1','0'),
            ('0','1','1','0','0','1','1','1','0','1','1','1','0','0'),
            ('0','1','1','0','0','1','1','1','0','1','1','1','1','0'),
            ('0','1','1','0','0','1','1','1','1','0','0','0','0','0'),
            ('0','1','1','0','0','1','1','1','1','0','0','0','1','0'),
            ('0','1','1','0','0','1','1','1','1','0','0','1','0','0'),
            ('0','1','1','0','0','1','1','1','1','0','0','1','1','0'),
            ('0','1','1','0','0','1','1','1','1','0','1','0','0','0'),
            ('0','1','1','0','0','1','1','1','1','0','1','0','1','0'),
            ('0','1','1','0','0','1','1','1','1','0','1','1','0','0'),
            ('0','1','1','0','0','1','1','1','1','0','1','1','1','0'),
            ('0','1','1','0','0','1','1','1','1','1','0','0','0','0'),
            ('0','1','1','0','0','1','1','1','1','1','0','0','1','0'),
            ('0','1','1','0','0','1','1','1','1','1','0','1','0','0'),
            ('0','1','1','0','0','1','1','1','1','1','0','1','1','0'),
            ('0','1','1','0','0','1','1','1','1','1','1','0','0','0'),
            ('0','1','1','0','0','1','1','1','1','1','1','0','1','0'),
            ('0','1','1','0','0','1','1','1','1','1','1','1','0','0'),
            ('0','1','1','0','0','1','1','1','1','1','1','1','1','0'),
            ('0','1','1','0','1','0','0','0','0','0','0','0','0','0'),
            ('0','1','1','0','1','0','0','0','0','0','0','0','1','0'),
            ('0','1','1','0','1','0','0','0','0','0','0','1','0','0'),
            ('0','1','1','0','1','0','0','0','0','0','0','1','1','0'),
            ('0','1','1','0','1','0','0','0','0','0','1','0','0','0'),
            ('0','1','1','0','1','0','0','0','0','0','1','0','1','0'),
            ('0','1','1','0','1','0','0','0','0','0','1','1','0','0'),
            ('0','1','1','0','1','0','0','0','0','0','1','1','1','0'),
            ('0','1','1','0','1','0','0','0','0','1','0','0','0','0'),
            ('0','1','1','0','1','0','0','0','0','1','0','0','1','0'),
            ('0','1','1','0','1','0','0','0','0','1','0','1','0','0'),
            ('0','1','1','0','1','0','0','0','0','1','0','1','1','0'),
            ('0','1','1','0','1','0','0','0','0','1','1','0','0','0'),
            ('0','1','1','0','1','0','0','0','0','1','1','0','1','0'),
            ('0','1','1','0','1','0','0','0','0','1','1','1','0','0'),
            ('0','1','1','0','1','0','0','0','0','1','1','1','1','0'),
            ('0','1','1','0','1','0','0','0','1','0','0','0','0','0'),
            ('0','1','1','0','1','0','0','0','1','0','0','0','1','0'),
            ('0','1','1','0','1','0','0','0','1','0','0','1','0','0'),
            ('0','1','1','0','1','0','0','0','1','0','0','1','1','0'),
            ('0','1','1','0','1','0','0','0','1','0','1','0','0','0'),
            ('0','1','1','0','1','0','0','0','1','0','1','0','1','0'),
            ('0','1','1','0','1','0','0','0','1','0','1','1','0','0'),
            ('0','1','1','0','1','0','0','0','1','0','1','1','1','0'),
            ('0','1','1','0','1','0','0','0','1','1','0','0','0','0'),
            ('0','1','1','0','1','0','0','0','1','1','0','0','1','0'),
            ('0','1','1','0','1','0','0','0','1','1','0','1','0','0'),
            ('0','1','1','0','1','0','0','0','1','1','0','1','1','0'),
            ('0','1','1','0','1','0','0','0','1','1','1','0','0','0'),
            ('0','1','1','0','1','0','0','0','1','1','1','0','1','0'),
            ('0','1','1','0','1','0','0','0','1','1','1','1','0','0'),
            ('0','1','1','0','1','0','0','0','1','1','1','1','1','0'),
            ('0','1','1','0','1','0','0','1','0','0','0','0','0','0'),
            ('0','1','1','0','1','0','0','1','0','0','0','0','1','0'),
            ('0','1','1','0','1','0','0','1','0','0','0','1','0','0'),
            ('0','1','1','0','1','0','0','1','0','0','0','1','1','0'),
            ('0','1','1','0','1','0','0','1','0','0','1','0','0','0'),
            ('0','1','1','0','1','0','0','1','0','0','1','0','1','0'),
            ('0','1','1','0','1','0','0','1','0','0','1','1','0','0'),
            ('0','1','1','0','1','0','0','1','0','0','1','1','1','0'),
            ('0','1','1','0','1','0','0','1','0','1','0','0','0','0'),
            ('0','1','1','0','1','0','0','1','0','1','0','0','1','0'),
            ('0','1','1','0','1','0','0','1','0','1','0','1','0','0'),
            ('0','1','1','0','1','0','0','1','0','1','0','1','1','0'),
            ('0','1','1','0','1','0','0','1','0','1','1','0','0','0'),
            ('0','1','1','0','1','0','0','1','0','1','1','0','1','0'),
            ('0','1','1','0','1','0','0','1','0','1','1','1','0','0'),
            ('0','1','1','0','1','0','0','1','0','1','1','1','1','0'),
            ('0','1','1','0','1','0','0','1','1','0','0','0','0','0'),
            ('0','1','1','0','1','0','0','1','1','0','0','0','1','0'),
            ('0','1','1','0','1','0','0','1','1','0','0','1','0','0'),
            ('0','1','1','0','1','0','0','1','1','0','0','1','1','0'),
            ('0','1','1','0','1','0','0','1','1','0','1','0','0','0'),
            ('0','1','1','0','1','0','0','1','1','0','1','0','1','0'),
            ('0','1','1','0','1','0','0','1','1','0','1','1','0','0'),
            ('0','1','1','0','1','0','0','1','1','0','1','1','1','0'),
            ('0','1','1','0','1','0','0','1','1','1','0','0','0','0'),
            ('0','1','1','0','1','0','0','1','1','1','0','0','1','0'),
            ('0','1','1','0','1','0','0','1','1','1','0','1','0','0'),
            ('0','1','1','0','1','0','0','1','1','1','0','1','1','0'),
            ('0','1','1','0','1','0','0','1','1','1','1','0','0','0'),
            ('0','1','1','0','1','0','0','1','1','1','1','0','1','0'),
            ('0','1','1','0','1','0','0','1','1','1','1','1','0','0'),
            ('0','1','1','0','1','0','0','1','1','1','1','1','1','0'),
            ('0','1','1','0','1','0','1','0','0','0','0','0','0','0'),
            ('0','1','1','0','1','0','1','0','0','0','0','0','1','0'),
            ('0','1','1','0','1','0','1','0','0','0','0','1','0','0'),
            ('0','1','1','0','1','0','1','0','0','0','0','1','1','0'),
            ('0','1','1','0','1','0','1','0','0','0','1','0','0','0'),
            ('0','1','1','0','1','0','1','0','0','0','1','0','1','0'),
            ('0','1','1','0','1','0','1','0','0','0','1','1','0','0'),
            ('0','1','1','0','1','0','1','0','0','0','1','1','1','0'),
            ('0','1','1','0','1','0','1','0','0','1','0','0','0','0'),
            ('0','1','1','0','1','0','1','0','0','1','0','0','1','0'),
            ('0','1','1','0','1','0','1','0','0','1','0','1','0','0'),
            ('0','1','1','0','1','0','1','0','0','1','0','1','1','0'),
            ('0','1','1','0','1','0','1','0','0','1','1','0','0','0'),
            ('0','1','1','0','1','0','1','0','0','1','1','0','1','0'),
            ('0','1','1','0','1','0','1','0','0','1','1','1','0','0'),
            ('0','1','1','0','1','0','1','0','0','1','1','1','1','0'),
            ('0','1','1','0','1','0','1','0','1','0','0','0','0','0'),
            ('0','1','1','0','1','0','1','0','1','0','0','0','1','0'),
            ('0','1','1','0','1','0','1','0','1','0','0','1','0','0'),
            ('0','1','1','0','1','0','1','0','1','0','0','1','1','0'),
            ('0','1','1','0','1','0','1','0','1','0','1','0','0','0'),
            ('0','1','1','0','1','0','1','0','1','0','1','0','1','0'),
            ('0','1','1','0','1','0','1','0','1','0','1','1','0','0'),
            ('0','1','1','0','1','0','1','0','1','0','1','1','1','0'),
            ('0','1','1','0','1','0','1','0','1','1','0','0','0','0'),
            ('0','1','1','0','1','0','1','0','1','1','0','0','1','0'),
            ('0','1','1','0','1','0','1','0','1','1','0','1','0','0'),
            ('0','1','1','0','1','0','1','0','1','1','0','1','1','0'),
            ('0','1','1','0','1','0','1','0','1','1','1','0','0','0'),
            ('0','1','1','0','1','0','1','0','1','1','1','0','1','0'),
            ('0','1','1','0','1','0','1','0','1','1','1','1','0','0'),
            ('0','1','1','0','1','0','1','0','1','1','1','1','1','0'),
            ('0','1','1','0','1','0','1','1','0','0','0','0','0','0'),
            ('0','1','1','0','1','0','1','1','0','0','0','0','1','0'),
            ('0','1','1','0','1','0','1','1','0','0','0','1','0','0'),
            ('0','1','1','0','1','0','1','1','0','0','0','1','1','0'),
            ('0','1','1','0','1','0','1','1','0','0','1','0','0','0'),
            ('0','1','1','0','1','0','1','1','0','0','1','0','1','0'),
            ('0','1','1','0','1','0','1','1','0','0','1','1','0','0'),
            ('0','1','1','0','1','0','1','1','0','0','1','1','1','0'),
            ('0','1','1','0','1','0','1','1','0','1','0','0','0','0'),
            ('0','1','1','0','1','0','1','1','0','1','0','0','1','0'),
            ('0','1','1','0','1','0','1','1','0','1','0','1','0','0'),
            ('0','1','1','0','1','0','1','1','0','1','0','1','1','0'),
            ('0','1','1','0','1','0','1','1','0','1','1','0','0','0'),
            ('0','1','1','0','1','0','1','1','0','1','1','0','1','0'),
            ('0','1','1','0','1','0','1','1','0','1','1','1','0','0'),
            ('0','1','1','0','1','0','1','1','0','1','1','1','1','0'),
            ('0','1','1','0','1','0','1','1','1','0','0','0','0','0'),
            ('0','1','1','0','1','0','1','1','1','0','0','0','1','0'),
            ('0','1','1','0','1','0','1','1','1','0','0','1','0','0'),
            ('0','1','1','0','1','0','1','1','1','0','0','1','1','0'),
            ('0','1','1','0','1','0','1','1','1','0','1','0','0','0'),
            ('0','1','1','0','1','0','1','1','1','0','1','0','1','0'),
            ('0','1','1','0','1','0','1','1','1','0','1','1','0','0'),
            ('0','1','1','0','1','0','1','1','1','0','1','1','1','0'),
            ('0','1','1','0','1','0','1','1','1','1','0','0','0','0'),
            ('0','1','1','0','1','0','1','1','1','1','0','0','1','0'),
            ('0','1','1','0','1','0','1','1','1','1','0','1','0','0'),
            ('0','1','1','0','1','0','1','1','1','1','0','1','1','0'),
            ('0','1','1','0','1','0','1','1','1','1','1','0','0','0'),
            ('0','1','1','0','1','0','1','1','1','1','1','0','1','0'),
            ('0','1','1','0','1','0','1','1','1','1','1','1','0','0'),
            ('0','1','1','0','1','0','1','1','1','1','1','1','1','0'),
            ('0','1','1','0','1','1','0','0','0','0','0','0','0','0'),
            ('0','1','1','0','1','1','0','0','0','0','0','0','1','0'),
            ('0','1','1','0','1','1','0','0','0','0','0','1','0','0'),
            ('0','1','1','0','1','1','0','0','0','0','0','1','1','0'),
            ('0','1','1','0','1','1','0','0','0','0','1','0','0','0'),
            ('0','1','1','0','1','1','0','0','0','0','1','0','1','0'),
            ('0','1','1','0','1','1','0','0','0','0','1','1','0','0'),
            ('0','1','1','0','1','1','0','0','0','0','1','1','1','0'),
            ('0','1','1','0','1','1','0','0','0','1','0','0','0','0'),
            ('0','1','1','0','1','1','0','0','0','1','0','0','1','0'),
            ('0','1','1','0','1','1','0','0','0','1','0','1','0','0'),
            ('0','1','1','0','1','1','0','0','0','1','0','1','1','0'),
            ('0','1','1','0','1','1','0','0','0','1','1','0','0','0'),
            ('0','1','1','0','1','1','0','0','0','1','1','0','1','0'),
            ('0','1','1','0','1','1','0','0','0','1','1','1','0','0'),
            ('0','1','1','0','1','1','0','0','0','1','1','1','1','0'),
            ('0','1','1','0','1','1','0','0','1','0','0','0','0','0'),
            ('0','1','1','0','1','1','0','0','1','0','0','0','1','0'),
            ('0','1','1','0','1','1','0','0','1','0','0','1','0','0'),
            ('0','1','1','0','1','1','0','0','1','0','0','1','1','0'),
            ('0','1','1','0','1','1','0','0','1','0','1','0','0','0'),
            ('0','1','1','0','1','1','0','0','1','0','1','0','1','0'),
            ('0','1','1','0','1','1','0','0','1','0','1','1','0','0'),
            ('0','1','1','0','1','1','0','0','1','0','1','1','1','0'),
            ('0','1','1','0','1','1','0','0','1','1','0','0','0','0'),
            ('0','1','1','0','1','1','0','0','1','1','0','0','1','0'),
            ('0','1','1','0','1','1','0','0','1','1','0','1','0','0'),
            ('0','1','1','0','1','1','0','0','1','1','0','1','1','0'),
            ('0','1','1','0','1','1','0','0','1','1','1','0','0','0'),
            ('0','1','1','0','1','1','0','0','1','1','1','0','1','0'),
            ('0','1','1','0','1','1','0','0','1','1','1','1','0','0'),
            ('0','1','1','0','1','1','0','0','1','1','1','1','1','0'),
            ('0','1','1','0','1','1','0','1','0','0','0','0','0','0'),
            ('0','1','1','0','1','1','0','1','0','0','0','0','1','0'),
            ('0','1','1','0','1','1','0','1','0','0','0','1','0','0'),
            ('0','1','1','0','1','1','0','1','0','0','0','1','1','0'),
            ('0','1','1','0','1','1','0','1','0','0','1','0','0','0'),
            ('0','1','1','0','1','1','0','1','0','0','1','0','1','0'),
            ('0','1','1','0','1','1','0','1','0','0','1','1','0','0'),
            ('0','1','1','0','1','1','0','1','0','0','1','1','1','0'),
            ('0','1','1','0','1','1','0','1','0','1','0','0','0','0'),
            ('0','1','1','0','1','1','0','1','0','1','0','0','1','0'),
            ('0','1','1','0','1','1','0','1','0','1','0','1','0','0'),
            ('0','1','1','0','1','1','0','1','0','1','0','1','1','0'),
            ('0','1','1','0','1','1','0','1','0','1','1','0','0','0'),
            ('0','1','1','0','1','1','0','1','0','1','1','0','1','0'),
            ('0','1','1','0','1','1','0','1','0','1','1','1','0','0'),
            ('0','1','1','0','1','1','0','1','0','1','1','1','1','0'),
            ('0','1','1','0','1','1','0','1','1','0','0','0','0','0'),
            ('0','1','1','0','1','1','0','1','1','0','0','0','1','0'),
            ('0','1','1','0','1','1','0','1','1','0','0','1','0','0'),
            ('0','1','1','0','1','1','0','1','1','0','0','1','1','0'),
            ('0','1','1','0','1','1','0','1','1','0','1','0','0','0'),
            ('0','1','1','0','1','1','0','1','1','0','1','0','1','0'),
            ('0','1','1','0','1','1','0','1','1','0','1','1','0','0'),
            ('0','1','1','0','1','1','0','1','1','0','1','1','1','0'),
            ('0','1','1','0','1','1','0','1','1','1','0','0','0','0'),
            ('0','1','1','0','1','1','0','1','1','1','0','0','1','0'),
            ('0','1','1','0','1','1','0','1','1','1','0','1','0','0'),
            ('0','1','1','0','1','1','0','1','1','1','0','1','1','0'),
            ('0','1','1','0','1','1','0','1','1','1','1','0','0','0'),
            ('0','1','1','0','1','1','0','1','1','1','1','0','1','0'),
            ('0','1','1','0','1','1','0','1','1','1','1','1','0','0'),
            ('0','1','1','0','1','1','0','1','1','1','1','1','1','0'),
            ('0','1','1','0','1','1','1','0','0','0','0','0','0','0'),
            ('0','1','1','0','1','1','1','0','0','0','0','0','1','0'),
            ('0','1','1','0','1','1','1','0','0','0','0','1','0','0'),
            ('0','1','1','0','1','1','1','0','0','0','0','1','1','0'),
            ('0','1','1','0','1','1','1','0','0','0','1','0','0','0'),
            ('0','1','1','0','1','1','1','0','0','0','1','0','1','0'),
            ('0','1','1','0','1','1','1','0','0','0','1','1','0','0'),
            ('0','1','1','0','1','1','1','0','0','0','1','1','1','0'),
            ('0','1','1','0','1','1','1','0','0','1','0','0','0','0'),
            ('0','1','1','0','1','1','1','0','0','1','0','0','1','0'),
            ('0','1','1','0','1','1','1','0','0','1','0','1','0','0'),
            ('0','1','1','0','1','1','1','0','0','1','0','1','1','0'),
            ('0','1','1','0','1','1','1','0','0','1','1','0','0','0'),
            ('0','1','1','0','1','1','1','0','0','1','1','0','1','0'),
            ('0','1','1','0','1','1','1','0','0','1','1','1','0','0'),
            ('0','1','1','0','1','1','1','0','0','1','1','1','1','0'),
            ('0','1','1','0','1','1','1','0','1','0','0','0','0','0'),
            ('0','1','1','0','1','1','1','0','1','0','0','0','1','0'),
            ('0','1','1','0','1','1','1','0','1','0','0','1','0','0'),
            ('0','1','1','0','1','1','1','0','1','0','0','1','1','0'),
            ('0','1','1','0','1','1','1','0','1','0','1','0','0','0'),
            ('0','1','1','0','1','1','1','0','1','0','1','0','1','0'),
            ('0','1','1','0','1','1','1','0','1','0','1','1','0','0'),
            ('0','1','1','0','1','1','1','0','1','0','1','1','1','0'),
            ('0','1','1','0','1','1','1','0','1','1','0','0','0','0'),
            ('0','1','1','0','1','1','1','0','1','1','0','0','1','0'),
            ('0','1','1','0','1','1','1','0','1','1','0','1','0','0'),
            ('0','1','1','0','1','1','1','0','1','1','0','1','1','0'),
            ('0','1','1','0','1','1','1','0','1','1','1','0','0','0'),
            ('0','1','1','0','1','1','1','0','1','1','1','0','1','0'),
            ('0','1','1','0','1','1','1','0','1','1','1','1','0','0'),
            ('0','1','1','0','1','1','1','0','1','1','1','1','1','0'),
            ('0','1','1','0','1','1','1','1','0','0','0','0','0','0'),
            ('0','1','1','0','1','1','1','1','0','0','0','0','1','0'),
            ('0','1','1','0','1','1','1','1','0','0','0','1','0','0'),
            ('0','1','1','0','1','1','1','1','0','0','0','1','1','0'),
            ('0','1','1','0','1','1','1','1','0','0','1','0','0','0'),
            ('0','1','1','0','1','1','1','1','0','0','1','0','1','0'),
            ('0','1','1','0','1','1','1','1','0','0','1','1','0','0'),
            ('0','1','1','0','1','1','1','1','0','0','1','1','1','0'),
            ('0','1','1','0','1','1','1','1','0','1','0','0','0','0'),
            ('0','1','1','0','1','1','1','1','0','1','0','0','1','0'),
            ('0','1','1','0','1','1','1','1','0','1','0','1','0','0'),
            ('0','1','1','0','1','1','1','1','0','1','0','1','1','0'),
            ('0','1','1','0','1','1','1','1','0','1','1','0','0','0'),
            ('0','1','1','0','1','1','1','1','0','1','1','0','1','0'),
            ('0','1','1','0','1','1','1','1','0','1','1','1','0','0'),
            ('0','1','1','0','1','1','1','1','0','1','1','1','1','0'),
            ('0','1','1','0','1','1','1','1','1','0','0','0','0','0'),
            ('0','1','1','0','1','1','1','1','1','0','0','0','1','0'),
            ('0','1','1','0','1','1','1','1','1','0','0','1','0','0'),
            ('0','1','1','0','1','1','1','1','1','0','0','1','1','0'),
            ('0','1','1','0','1','1','1','1','1','0','1','0','0','0'),
            ('0','1','1','0','1','1','1','1','1','0','1','0','1','0'),
            ('0','1','1','0','1','1','1','1','1','0','1','1','0','0'),
            ('0','1','1','0','1','1','1','1','1','0','1','1','1','0'),
            ('0','1','1','0','1','1','1','1','1','1','0','0','0','0'),
            ('0','1','1','0','1','1','1','1','1','1','0','0','1','0'),
            ('0','1','1','0','1','1','1','1','1','1','0','1','0','0'),
            ('0','1','1','0','1','1','1','1','1','1','0','1','1','0'),
            ('0','1','1','0','1','1','1','1','1','1','1','0','0','0'),
            ('0','1','1','0','1','1','1','1','1','1','1','0','1','0'),
            ('0','1','1','0','1','1','1','1','1','1','1','1','0','0'),
            ('0','1','1','0','1','1','1','1','1','1','1','1','1','0'),
            ('0','1','1','1','0','0','0','0','0','0','0','0','0','0'),
            ('0','1','1','1','0','0','0','0','0','0','0','0','1','0'),
            ('0','1','1','1','0','0','0','0','0','0','0','1','0','0'),
            ('0','1','1','1','0','0','0','0','0','0','0','1','1','0'),
            ('0','1','1','1','0','0','0','0','0','0','1','0','0','0'),
            ('0','1','1','1','0','0','0','0','0','0','1','0','1','0'),
            ('0','1','1','1','0','0','0','0','0','0','1','1','0','0'),
            ('0','1','1','1','0','0','0','0','0','0','1','1','1','0'),
            ('0','1','1','1','0','0','0','0','0','1','0','0','0','0'),
            ('0','1','1','1','0','0','0','0','0','1','0','0','1','0'),
            ('0','1','1','1','0','0','0','0','0','1','0','1','0','0'),
            ('0','1','1','1','0','0','0','0','0','1','0','1','1','0'),
            ('0','1','1','1','0','0','0','0','0','1','1','0','0','0'),
            ('0','1','1','1','0','0','0','0','0','1','1','0','1','0'),
            ('0','1','1','1','0','0','0','0','0','1','1','1','0','0'),
            ('0','1','1','1','0','0','0','0','0','1','1','1','1','0'),
            ('0','1','1','1','0','0','0','0','1','0','0','0','0','0'),
            ('0','1','1','1','0','0','0','0','1','0','0','0','1','0'),
            ('0','1','1','1','0','0','0','0','1','0','0','1','0','0'),
            ('0','1','1','1','0','0','0','0','1','0','0','1','1','0'),
            ('0','1','1','1','0','0','0','0','1','0','1','0','0','0'),
            ('0','1','1','1','0','0','0','0','1','0','1','0','1','0'),
            ('0','1','1','1','0','0','0','0','1','0','1','1','0','0'),
            ('0','1','1','1','0','0','0','0','1','0','1','1','1','0'),
            ('0','1','1','1','0','0','0','0','1','1','0','0','0','0'),
            ('0','1','1','1','0','0','0','0','1','1','0','0','1','0'),
            ('0','1','1','1','0','0','0','0','1','1','0','1','0','0'),
            ('0','1','1','1','0','0','0','0','1','1','0','1','1','0'),
            ('0','1','1','1','0','0','0','0','1','1','1','0','0','0'),
            ('0','1','1','1','0','0','0','0','1','1','1','0','1','0'),
            ('0','1','1','1','0','0','0','0','1','1','1','1','0','0'),
            ('0','1','1','1','0','0','0','0','1','1','1','1','1','0'),
            ('0','1','1','1','0','0','0','1','0','0','0','0','0','0'),
            ('0','1','1','1','0','0','0','1','0','0','0','0','1','0'),
            ('0','1','1','1','0','0','0','1','0','0','0','1','0','0'),
            ('0','1','1','1','0','0','0','1','0','0','0','1','1','0'),
            ('0','1','1','1','0','0','0','1','0','0','1','0','0','0'),
            ('0','1','1','1','0','0','0','1','0','0','1','0','1','0'),
            ('0','1','1','1','0','0','0','1','0','0','1','1','0','0'),
            ('0','1','1','1','0','0','0','1','0','0','1','1','1','0'),
            ('0','1','1','1','0','0','0','1','0','1','0','0','0','0'),
            ('0','1','1','1','0','0','0','1','0','1','0','0','1','0'),
            ('0','1','1','1','0','0','0','1','0','1','0','1','0','0'),
            ('0','1','1','1','0','0','0','1','0','1','0','1','1','0'),
            ('0','1','1','1','0','0','0','1','0','1','1','0','0','0'),
            ('0','1','1','1','0','0','0','1','0','1','1','0','1','0'),
            ('0','1','1','1','0','0','0','1','0','1','1','1','0','0'),
            ('0','1','1','1','0','0','0','1','0','1','1','1','1','0'),
            ('0','1','1','1','0','0','0','1','1','0','0','0','0','0'),
            ('0','1','1','1','0','0','0','1','1','0','0','0','1','0'),
            ('0','1','1','1','0','0','0','1','1','0','0','1','0','0'),
            ('0','1','1','1','0','0','0','1','1','0','0','1','1','0'),
            ('0','1','1','1','0','0','0','1','1','0','1','0','0','0'),
            ('0','1','1','1','0','0','0','1','1','0','1','0','1','0'),
            ('0','1','1','1','0','0','0','1','1','0','1','1','0','0'),
            ('0','1','1','1','0','0','0','1','1','0','1','1','1','0'),
            ('0','1','1','1','0','0','0','1','1','1','0','0','0','0'),
            ('0','1','1','1','0','0','0','1','1','1','0','0','1','0'),
            ('0','1','1','1','0','0','0','1','1','1','0','1','0','0'),
            ('0','1','1','1','0','0','0','1','1','1','0','1','1','0'),
            ('0','1','1','1','0','0','0','1','1','1','1','0','0','0'),
            ('0','1','1','1','0','0','0','1','1','1','1','0','1','0'),
            ('0','1','1','1','0','0','0','1','1','1','1','1','0','0'),
            ('0','1','1','1','0','0','0','1','1','1','1','1','1','0'),
            ('0','1','1','1','0','0','1','0','0','0','0','0','0','0'),
            ('0','1','1','1','0','0','1','0','0','0','0','0','1','0'),
            ('0','1','1','1','0','0','1','0','0','0','0','1','0','0'),
            ('0','1','1','1','0','0','1','0','0','0','0','1','1','0'),
            ('0','1','1','1','0','0','1','0','0','0','1','0','0','0'),
            ('0','1','1','1','0','0','1','0','0','0','1','0','1','0'),
            ('0','1','1','1','0','0','1','0','0','0','1','1','0','0'),
            ('0','1','1','1','0','0','1','0','0','0','1','1','1','0'),
            ('0','1','1','1','0','0','1','0','0','1','0','0','0','0'),
            ('0','1','1','1','0','0','1','0','0','1','0','0','1','0'),
            ('0','1','1','1','0','0','1','0','0','1','0','1','0','0'),
            ('0','1','1','1','0','0','1','0','0','1','0','1','1','0'),
            ('0','1','1','1','0','0','1','0','0','1','1','0','0','0'),
            ('0','1','1','1','0','0','1','0','0','1','1','0','1','0'),
            ('0','1','1','1','0','0','1','0','0','1','1','1','0','0'),
            ('0','1','1','1','0','0','1','0','0','1','1','1','1','0'),
            ('0','1','1','1','0','0','1','0','1','0','0','0','0','0'),
            ('0','1','1','1','0','0','1','0','1','0','0','0','1','0'),
            ('0','1','1','1','0','0','1','0','1','0','0','1','0','0'),
            ('0','1','1','1','0','0','1','0','1','0','0','1','1','0'),
            ('0','1','1','1','0','0','1','0','1','0','1','0','0','0'),
            ('0','1','1','1','0','0','1','0','1','0','1','0','1','0'),
            ('0','1','1','1','0','0','1','0','1','0','1','1','0','0'),
            ('0','1','1','1','0','0','1','0','1','0','1','1','1','0'),
            ('0','1','1','1','0','0','1','0','1','1','0','0','0','0'),
            ('0','1','1','1','0','0','1','0','1','1','0','0','1','0'),
            ('0','1','1','1','0','0','1','0','1','1','0','1','0','0'),
            ('0','1','1','1','0','0','1','0','1','1','0','1','1','0'),
            ('0','1','1','1','0','0','1','0','1','1','1','0','0','0'),
            ('0','1','1','1','0','0','1','0','1','1','1','0','1','0'),
            ('0','1','1','1','0','0','1','0','1','1','1','1','0','0'),
            ('0','1','1','1','0','0','1','0','1','1','1','1','1','0'),
            ('0','1','1','1','0','0','1','1','0','0','0','0','0','0'),
            ('0','1','1','1','0','0','1','1','0','0','0','0','1','0'),
            ('0','1','1','1','0','0','1','1','0','0','0','1','0','0'),
            ('0','1','1','1','0','0','1','1','0','0','0','1','1','0'),
            ('0','1','1','1','0','0','1','1','0','0','1','0','0','0'),
            ('0','1','1','1','0','0','1','1','0','0','1','0','1','0'),
            ('0','1','1','1','0','0','1','1','0','0','1','1','0','0'),
            ('0','1','1','1','0','0','1','1','0','0','1','1','1','0'),
            ('0','1','1','1','0','0','1','1','0','1','0','0','0','0'),
            ('0','1','1','1','0','0','1','1','0','1','0','0','1','0'),
            ('0','1','1','1','0','0','1','1','0','1','0','1','0','0'),
            ('0','1','1','1','0','0','1','1','0','1','0','1','1','0'),
            ('0','1','1','1','0','0','1','1','0','1','1','0','0','0'),
            ('0','1','1','1','0','0','1','1','0','1','1','0','1','0'),
            ('0','1','1','1','0','0','1','1','0','1','1','1','0','0'),
            ('0','1','1','1','0','0','1','1','0','1','1','1','1','0'),
            ('0','1','1','1','0','0','1','1','1','0','0','0','0','0'),
            ('0','1','1','1','0','0','1','1','1','0','0','0','1','0'),
            ('0','1','1','1','0','0','1','1','1','0','0','1','0','0'),
            ('0','1','1','1','0','0','1','1','1','0','0','1','1','0'),
            ('0','1','1','1','0','0','1','1','1','0','1','0','0','0'),
            ('0','1','1','1','0','0','1','1','1','0','1','0','1','0'),
            ('0','1','1','1','0','0','1','1','1','0','1','1','0','0'),
            ('0','1','1','1','0','0','1','1','1','0','1','1','1','0'),
            ('0','1','1','1','0','0','1','1','1','1','0','0','0','0'),
            ('0','1','1','1','0','0','1','1','1','1','0','0','1','0'),
            ('0','1','1','1','0','0','1','1','1','1','0','1','0','0'),
            ('0','1','1','1','0','0','1','1','1','1','0','1','1','0'),
            ('0','1','1','1','0','0','1','1','1','1','1','0','0','0'),
            ('0','1','1','1','0','0','1','1','1','1','1','0','1','0'),
            ('0','1','1','1','0','0','1','1','1','1','1','1','0','0'),
            ('0','1','1','1','0','0','1','1','1','1','1','1','1','0'),
            ('0','1','1','1','0','1','0','0','0','0','0','0','0','0'),
            ('0','1','1','1','0','1','0','0','0','0','0','0','1','0'),
            ('0','1','1','1','0','1','0','0','0','0','0','1','0','0'),
            ('0','1','1','1','0','1','0','0','0','0','0','1','1','0'),
            ('0','1','1','1','0','1','0','0','0','0','1','0','0','0'),
            ('0','1','1','1','0','1','0','0','0','0','1','0','1','0'),
            ('0','1','1','1','0','1','0','0','0','0','1','1','0','0'),
            ('0','1','1','1','0','1','0','0','0','0','1','1','1','0'),
            ('0','1','1','1','0','1','0','0','0','1','0','0','0','0'),
            ('0','1','1','1','0','1','0','0','0','1','0','0','1','0'),
            ('0','1','1','1','0','1','0','0','0','1','0','1','0','0'),
            ('0','1','1','1','0','1','0','0','0','1','0','1','1','0'),
            ('0','1','1','1','0','1','0','0','0','1','1','0','0','0'),
            ('0','1','1','1','0','1','0','0','0','1','1','0','1','0'),
            ('0','1','1','1','0','1','0','0','0','1','1','1','0','0'),
            ('0','1','1','1','0','1','0','0','0','1','1','1','1','0'),
            ('0','1','1','1','0','1','0','0','1','0','0','0','0','0'),
            ('0','1','1','1','0','1','0','0','1','0','0','0','1','0'),
            ('0','1','1','1','0','1','0','0','1','0','0','1','0','0'),
            ('0','1','1','1','0','1','0','0','1','0','0','1','1','0'),
            ('0','1','1','1','0','1','0','0','1','0','1','0','0','0'),
            ('0','1','1','1','0','1','0','0','1','0','1','0','1','0'),
            ('0','1','1','1','0','1','0','0','1','0','1','1','0','0'),
            ('0','1','1','1','0','1','0','0','1','0','1','1','1','0'),
            ('0','1','1','1','0','1','0','0','1','1','0','0','0','0'),
            ('0','1','1','1','0','1','0','0','1','1','0','0','1','0'),
            ('0','1','1','1','0','1','0','0','1','1','0','1','0','0'),
            ('0','1','1','1','0','1','0','0','1','1','0','1','1','0'),
            ('0','1','1','1','0','1','0','0','1','1','1','0','0','0'),
            ('0','1','1','1','0','1','0','0','1','1','1','0','1','0'),
            ('0','1','1','1','0','1','0','0','1','1','1','1','0','0'),
            ('0','1','1','1','0','1','0','0','1','1','1','1','1','0'),
            ('0','1','1','1','0','1','0','1','0','0','0','0','0','0'),
            ('0','1','1','1','0','1','0','1','0','0','0','0','1','0'),
            ('0','1','1','1','0','1','0','1','0','0','0','1','0','0'),
            ('0','1','1','1','0','1','0','1','0','0','0','1','1','0'),
            ('0','1','1','1','0','1','0','1','0','0','1','0','0','0'),
            ('0','1','1','1','0','1','0','1','0','0','1','0','1','0'),
            ('0','1','1','1','0','1','0','1','0','0','1','1','0','0'),
            ('0','1','1','1','0','1','0','1','0','0','1','1','1','0'),
            ('0','1','1','1','0','1','0','1','0','1','0','0','0','0'),
            ('0','1','1','1','0','1','0','1','0','1','0','0','1','0'),
            ('0','1','1','1','0','1','0','1','0','1','0','1','0','0'),
            ('0','1','1','1','0','1','0','1','0','1','0','1','1','0'),
            ('0','1','1','1','0','1','0','1','0','1','1','0','0','0'),
            ('0','1','1','1','0','1','0','1','0','1','1','0','1','0'),
            ('0','1','1','1','0','1','0','1','0','1','1','1','0','0'),
            ('0','1','1','1','0','1','0','1','0','1','1','1','1','0'),
            ('0','1','1','1','0','1','0','1','1','0','0','0','0','0'),
            ('0','1','1','1','0','1','0','1','1','0','0','0','1','0'),
            ('0','1','1','1','0','1','0','1','1','0','0','1','0','0'),
            ('0','1','1','1','0','1','0','1','1','0','0','1','1','0'),
            ('0','1','1','1','0','1','0','1','1','0','1','0','0','0'),
            ('0','1','1','1','0','1','0','1','1','0','1','0','1','0'),
            ('0','1','1','1','0','1','0','1','1','0','1','1','0','0'),
            ('0','1','1','1','0','1','0','1','1','0','1','1','1','0'),
            ('0','1','1','1','0','1','0','1','1','1','0','0','0','0'),
            ('0','1','1','1','0','1','0','1','1','1','0','0','1','0'),
            ('0','1','1','1','0','1','0','1','1','1','0','1','0','0'),
            ('0','1','1','1','0','1','0','1','1','1','0','1','1','0'),
            ('0','1','1','1','0','1','0','1','1','1','1','0','0','0'),
            ('0','1','1','1','0','1','0','1','1','1','1','0','1','0'),
            ('0','1','1','1','0','1','0','1','1','1','1','1','0','0'),
            ('0','1','1','1','0','1','0','1','1','1','1','1','1','0'),
            ('0','1','1','1','0','1','1','0','0','0','0','0','0','0'),
            ('0','1','1','1','0','1','1','0','0','0','0','0','1','0'),
            ('0','1','1','1','0','1','1','0','0','0','0','1','0','0'),
            ('0','1','1','1','0','1','1','0','0','0','0','1','1','0'),
            ('0','1','1','1','0','1','1','0','0','0','1','0','0','0'),
            ('0','1','1','1','0','1','1','0','0','0','1','0','1','0'),
            ('0','1','1','1','0','1','1','0','0','0','1','1','0','0'),
            ('0','1','1','1','0','1','1','0','0','0','1','1','1','0'),
            ('0','1','1','1','0','1','1','0','0','1','0','0','0','0'),
            ('0','1','1','1','0','1','1','0','0','1','0','0','1','0'),
            ('0','1','1','1','0','1','1','0','0','1','0','1','0','0'),
            ('0','1','1','1','0','1','1','0','0','1','0','1','1','0'),
            ('0','1','1','1','0','1','1','0','0','1','1','0','0','0'),
            ('0','1','1','1','0','1','1','0','0','1','1','0','1','0'),
            ('0','1','1','1','0','1','1','0','0','1','1','1','0','0'),
            ('0','1','1','1','0','1','1','0','0','1','1','1','1','0'),
            ('0','1','1','1','0','1','1','0','1','0','0','0','0','0'),
            ('0','1','1','1','0','1','1','0','1','0','0','0','1','0'),
            ('0','1','1','1','0','1','1','0','1','0','0','1','0','0'),
            ('0','1','1','1','0','1','1','0','1','0','0','1','1','0'),
            ('0','1','1','1','0','1','1','0','1','0','1','0','0','0'),
            ('0','1','1','1','0','1','1','0','1','0','1','0','1','0'),
            ('0','1','1','1','0','1','1','0','1','0','1','1','0','0'),
            ('0','1','1','1','0','1','1','0','1','0','1','1','1','0'),
            ('0','1','1','1','0','1','1','0','1','1','0','0','0','0'),
            ('0','1','1','1','0','1','1','0','1','1','0','0','1','0'),
            ('0','1','1','1','0','1','1','0','1','1','0','1','0','0'),
            ('0','1','1','1','0','1','1','0','1','1','0','1','1','0'),
            ('0','1','1','1','0','1','1','0','1','1','1','0','0','0'),
            ('0','1','1','1','0','1','1','0','1','1','1','0','1','0'),
            ('0','1','1','1','0','1','1','0','1','1','1','1','0','0'),
            ('0','1','1','1','0','1','1','0','1','1','1','1','1','0'),
            ('0','1','1','1','0','1','1','1','0','0','0','0','0','0'),
            ('0','1','1','1','0','1','1','1','0','0','0','0','1','0'),
            ('0','1','1','1','0','1','1','1','0','0','0','1','0','0'),
            ('0','1','1','1','0','1','1','1','0','0','0','1','1','0'),
            ('0','1','1','1','0','1','1','1','0','0','1','0','0','0'),
            ('0','1','1','1','0','1','1','1','0','0','1','0','1','0'),
            ('0','1','1','1','0','1','1','1','0','0','1','1','0','0'),
            ('0','1','1','1','0','1','1','1','0','0','1','1','1','0'),
            ('0','1','1','1','0','1','1','1','0','1','0','0','0','0'),
            ('0','1','1','1','0','1','1','1','0','1','0','0','1','0'),
            ('0','1','1','1','0','1','1','1','0','1','0','1','0','0'),
            ('0','1','1','1','0','1','1','1','0','1','0','1','1','0'),
            ('0','1','1','1','0','1','1','1','0','1','1','0','0','0'),
            ('0','1','1','1','0','1','1','1','0','1','1','0','1','0'),
            ('0','1','1','1','0','1','1','1','0','1','1','1','0','0'),
            ('0','1','1','1','0','1','1','1','0','1','1','1','1','0'),
            ('0','1','1','1','0','1','1','1','1','0','0','0','0','0'),
            ('0','1','1','1','0','1','1','1','1','0','0','0','1','0'),
            ('0','1','1','1','0','1','1','1','1','0','0','1','0','0'),
            ('0','1','1','1','0','1','1','1','1','0','0','1','1','0'),
            ('0','1','1','1','0','1','1','1','1','0','1','0','0','0'),
            ('0','1','1','1','0','1','1','1','1','0','1','0','1','0'),
            ('0','1','1','1','0','1','1','1','1','0','1','1','0','0'),
            ('0','1','1','1','0','1','1','1','1','0','1','1','1','0'),
            ('0','1','1','1','0','1','1','1','1','1','0','0','0','0'),
            ('0','1','1','1','0','1','1','1','1','1','0','0','1','0'),
            ('0','1','1','1','0','1','1','1','1','1','0','1','0','0'),
            ('0','1','1','1','0','1','1','1','1','1','0','1','1','0'),
            ('0','1','1','1','0','1','1','1','1','1','1','0','0','0'),
            ('0','1','1','1','0','1','1','1','1','1','1','0','1','0'),
            ('0','1','1','1','0','1','1','1','1','1','1','1','0','0'),
            ('0','1','1','1','0','1','1','1','1','1','1','1','1','0'),
            ('0','1','1','1','1','0','0','0','0','0','0','0','0','0'),
            ('0','1','1','1','1','0','0','0','0','0','0','0','1','0'),
            ('0','1','1','1','1','0','0','0','0','0','0','1','0','0'),
            ('0','1','1','1','1','0','0','0','0','0','0','1','1','0'),
            ('0','1','1','1','1','0','0','0','0','0','1','0','0','0'),
            ('0','1','1','1','1','0','0','0','0','0','1','0','1','0'),
            ('0','1','1','1','1','0','0','0','0','0','1','1','0','0'),
            ('0','1','1','1','1','0','0','0','0','0','1','1','1','0'),
            ('0','1','1','1','1','0','0','0','0','1','0','0','0','0'),
            ('0','1','1','1','1','0','0','0','0','1','0','0','1','0'),
            ('0','1','1','1','1','0','0','0','0','1','0','1','0','0'),
            ('0','1','1','1','1','0','0','0','0','1','0','1','1','0'),
            ('0','1','1','1','1','0','0','0','0','1','1','0','0','0'),
            ('0','1','1','1','1','0','0','0','0','1','1','0','1','0'),
            ('0','1','1','1','1','0','0','0','0','1','1','1','0','0'),
            ('0','1','1','1','1','0','0','0','0','1','1','1','1','0'),
            ('0','1','1','1','1','0','0','0','1','0','0','0','0','0'),
            ('0','1','1','1','1','0','0','0','1','0','0','0','1','0'),
            ('0','1','1','1','1','0','0','0','1','0','0','1','0','0'),
            ('0','1','1','1','1','0','0','0','1','0','0','1','1','0'),
            ('0','1','1','1','1','0','0','0','1','0','1','0','0','0'),
            ('0','1','1','1','1','0','0','0','1','0','1','0','1','0'),
            ('0','1','1','1','1','0','0','0','1','0','1','1','0','0'),
            ('0','1','1','1','1','0','0','0','1','0','1','1','1','0'),
            ('0','1','1','1','1','0','0','0','1','1','0','0','0','0'),
            ('0','1','1','1','1','0','0','0','1','1','0','0','1','0'),
            ('0','1','1','1','1','0','0','0','1','1','0','1','0','0'),
            ('0','1','1','1','1','0','0','0','1','1','0','1','1','0'),
            ('0','1','1','1','1','0','0','0','1','1','1','0','0','0'),
            ('0','1','1','1','1','0','0','0','1','1','1','0','1','0'),
            ('0','1','1','1','1','0','0','0','1','1','1','1','0','0'),
            ('0','1','1','1','1','0','0','0','1','1','1','1','1','0'),
            ('0','1','1','1','1','0','0','1','0','0','0','0','0','0'),
            ('0','1','1','1','1','0','0','1','0','0','0','0','1','0'),
            ('0','1','1','1','1','0','0','1','0','0','0','1','0','0'),
            ('0','1','1','1','1','0','0','1','0','0','0','1','1','0'),
            ('0','1','1','1','1','0','0','1','0','0','1','0','0','0'),
            ('0','1','1','1','1','0','0','1','0','0','1','0','1','0'),
            ('0','1','1','1','1','0','0','1','0','0','1','1','0','0'),
            ('0','1','1','1','1','0','0','1','0','0','1','1','1','0'),
            ('0','1','1','1','1','0','0','1','0','1','0','0','0','0'),
            ('0','1','1','1','1','0','0','1','0','1','0','0','1','0'),
            ('0','1','1','1','1','0','0','1','0','1','0','1','0','0'),
            ('0','1','1','1','1','0','0','1','0','1','0','1','1','0'),
            ('0','1','1','1','1','0','0','1','0','1','1','0','0','0'),
            ('0','1','1','1','1','0','0','1','0','1','1','0','1','0'),
            ('0','1','1','1','1','0','0','1','0','1','1','1','0','0'),
            ('0','1','1','1','1','0','0','1','0','1','1','1','1','0'),
            ('0','1','1','1','1','0','0','1','1','0','0','0','0','0'),
            ('0','1','1','1','1','0','0','1','1','0','0','0','1','0'),
            ('0','1','1','1','1','0','0','1','1','0','0','1','0','0'),
            ('0','1','1','1','1','0','0','1','1','0','0','1','1','0'),
            ('0','1','1','1','1','0','0','1','1','0','1','0','0','0'),
            ('0','1','1','1','1','0','0','1','1','0','1','0','1','0'),
            ('0','1','1','1','1','0','0','1','1','0','1','1','0','0'),
            ('0','1','1','1','1','0','0','1','1','0','1','1','1','0'),
            ('0','1','1','1','1','0','0','1','1','1','0','0','0','0'),
            ('0','1','1','1','1','0','0','1','1','1','0','0','1','0'),
            ('0','1','1','1','1','0','0','1','1','1','0','1','0','0'),
            ('0','1','1','1','1','0','0','1','1','1','0','1','1','0'),
            ('0','1','1','1','1','0','0','1','1','1','1','0','0','0'),
            ('0','1','1','1','1','0','0','1','1','1','1','0','1','0'),
            ('0','1','1','1','1','0','0','1','1','1','1','1','0','0'),
            ('0','1','1','1','1','0','0','1','1','1','1','1','1','0'),
            ('0','1','1','1','1','0','1','0','0','0','0','0','0','0'),
            ('0','1','1','1','1','0','1','0','0','0','0','0','1','0'),
            ('0','1','1','1','1','0','1','0','0','0','0','1','0','0'),
            ('0','1','1','1','1','0','1','0','0','0','0','1','1','0'),
            ('0','1','1','1','1','0','1','0','0','0','1','0','0','0'),
            ('0','1','1','1','1','0','1','0','0','0','1','0','1','0'),
            ('0','1','1','1','1','0','1','0','0','0','1','1','0','0'),
            ('0','1','1','1','1','0','1','0','0','0','1','1','1','0'),
            ('0','1','1','1','1','0','1','0','0','1','0','0','0','0'),
            ('0','1','1','1','1','0','1','0','0','1','0','0','1','0'),
            ('0','1','1','1','1','0','1','0','0','1','0','1','0','0'),
            ('0','1','1','1','1','0','1','0','0','1','0','1','1','0'),
            ('0','1','1','1','1','0','1','0','0','1','1','0','0','0'),
            ('0','1','1','1','1','0','1','0','0','1','1','0','1','0'),
            ('0','1','1','1','1','0','1','0','0','1','1','1','0','0'),
            ('0','1','1','1','1','0','1','0','0','1','1','1','1','0'),
            ('0','1','1','1','1','0','1','0','1','0','0','0','0','0'),
            ('0','1','1','1','1','0','1','0','1','0','0','0','1','0'),
            ('0','1','1','1','1','0','1','0','1','0','0','1','0','0'),
            ('0','1','1','1','1','0','1','0','1','0','0','1','1','0'),
            ('0','1','1','1','1','0','1','0','1','0','1','0','0','0'),
            ('0','1','1','1','1','0','1','0','1','0','1','0','1','0'),
            ('0','1','1','1','1','0','1','0','1','0','1','1','0','0'),
            ('0','1','1','1','1','0','1','0','1','0','1','1','1','0'),
            ('0','1','1','1','1','0','1','0','1','1','0','0','0','0'),
            ('0','1','1','1','1','0','1','0','1','1','0','0','1','0'),
            ('0','1','1','1','1','0','1','0','1','1','0','1','0','0'),
            ('0','1','1','1','1','0','1','0','1','1','0','1','1','0'),
            ('0','1','1','1','1','0','1','0','1','1','1','0','0','0'),
            ('0','1','1','1','1','0','1','0','1','1','1','0','1','0'),
            ('0','1','1','1','1','0','1','0','1','1','1','1','0','0'),
            ('0','1','1','1','1','0','1','0','1','1','1','1','1','0'),
            ('0','1','1','1','1','0','1','1','0','0','0','0','0','0'),
            ('0','1','1','1','1','0','1','1','0','0','0','0','1','0'),
            ('0','1','1','1','1','0','1','1','0','0','0','1','0','0'),
            ('0','1','1','1','1','0','1','1','0','0','0','1','1','0'),
            ('0','1','1','1','1','0','1','1','0','0','1','0','0','0'),
            ('0','1','1','1','1','0','1','1','0','0','1','0','1','0'),
            ('0','1','1','1','1','0','1','1','0','0','1','1','0','0'),
            ('0','1','1','1','1','0','1','1','0','0','1','1','1','0'),
            ('0','1','1','1','1','0','1','1','0','1','0','0','0','0'),
            ('0','1','1','1','1','0','1','1','0','1','0','0','1','0'),
            ('0','1','1','1','1','0','1','1','0','1','0','1','0','0'),
            ('0','1','1','1','1','0','1','1','0','1','0','1','1','0'),
            ('0','1','1','1','1','0','1','1','0','1','1','0','0','0'),
            ('0','1','1','1','1','0','1','1','0','1','1','0','1','0'),
            ('0','1','1','1','1','0','1','1','0','1','1','1','0','0'),
            ('0','1','1','1','1','0','1','1','0','1','1','1','1','0'),
            ('0','1','1','1','1','0','1','1','1','0','0','0','0','0'),
            ('0','1','1','1','1','0','1','1','1','0','0','0','1','0'),
            ('0','1','1','1','1','0','1','1','1','0','0','1','0','0'),
            ('0','1','1','1','1','0','1','1','1','0','0','1','1','0'),
            ('0','1','1','1','1','0','1','1','1','0','1','0','0','0'),
            ('0','1','1','1','1','0','1','1','1','0','1','0','1','0'),
            ('0','1','1','1','1','0','1','1','1','0','1','1','0','0'),
            ('0','1','1','1','1','0','1','1','1','0','1','1','1','0'),
            ('0','1','1','1','1','0','1','1','1','1','0','0','0','0'),
            ('0','1','1','1','1','0','1','1','1','1','0','0','1','0'),
            ('0','1','1','1','1','0','1','1','1','1','0','1','0','0'),
            ('0','1','1','1','1','0','1','1','1','1','0','1','1','0'),
            ('0','1','1','1','1','0','1','1','1','1','1','0','0','0'),
            ('0','1','1','1','1','0','1','1','1','1','1','0','1','0'),
            ('0','1','1','1','1','0','1','1','1','1','1','1','0','0'),
            ('0','1','1','1','1','0','1','1','1','1','1','1','1','0'),
            ('0','1','1','1','1','1','0','0','0','0','0','0','0','0'),
            ('0','1','1','1','1','1','0','0','0','0','0','0','1','0'),
            ('0','1','1','1','1','1','0','0','0','0','0','1','0','0'),
            ('0','1','1','1','1','1','0','0','0','0','0','1','1','0'),
            ('0','1','1','1','1','1','0','0','0','0','1','0','0','0'),
            ('0','1','1','1','1','1','0','0','0','0','1','0','1','0'),
            ('0','1','1','1','1','1','0','0','0','0','1','1','0','0'),
            ('0','1','1','1','1','1','0','0','0','0','1','1','1','0'),
            ('0','1','1','1','1','1','0','0','0','1','0','0','0','0'),
            ('0','1','1','1','1','1','0','0','0','1','0','0','1','0'),
            ('0','1','1','1','1','1','0','0','0','1','0','1','0','0'),
            ('0','1','1','1','1','1','0','0','0','1','0','1','1','0'),
            ('0','1','1','1','1','1','0','0','0','1','1','0','0','0'),
            ('0','1','1','1','1','1','0','0','0','1','1','0','1','0'),
            ('0','1','1','1','1','1','0','0','0','1','1','1','0','0'),
            ('0','1','1','1','1','1','0','0','0','1','1','1','1','0'),
            ('0','1','1','1','1','1','0','0','1','0','0','0','0','0'),
            ('0','1','1','1','1','1','0','0','1','0','0','0','1','0'),
            ('0','1','1','1','1','1','0','0','1','0','0','1','0','0'),
            ('0','1','1','1','1','1','0','0','1','0','0','1','1','0'),
            ('0','1','1','1','1','1','0','0','1','0','1','0','0','0'),
            ('0','1','1','1','1','1','0','0','1','0','1','0','1','0'),
            ('0','1','1','1','1','1','0','0','1','0','1','1','0','0'),
            ('0','1','1','1','1','1','0','0','1','0','1','1','1','0'),
            ('0','1','1','1','1','1','0','0','1','1','0','0','0','0'),
            ('0','1','1','1','1','1','0','0','1','1','0','0','1','0'),
            ('0','1','1','1','1','1','0','0','1','1','0','1','0','0'),
            ('0','1','1','1','1','1','0','0','1','1','0','1','1','0'),
            ('0','1','1','1','1','1','0','0','1','1','1','0','0','0'),
            ('0','1','1','1','1','1','0','0','1','1','1','0','1','0'),
            ('0','1','1','1','1','1','0','0','1','1','1','1','0','0'),
            ('0','1','1','1','1','1','0','0','1','1','1','1','1','0'),
            ('0','1','1','1','1','1','0','1','0','0','0','0','0','0'),
            ('0','1','1','1','1','1','0','1','0','0','0','0','1','0'),
            ('0','1','1','1','1','1','0','1','0','0','0','1','0','0'),
            ('0','1','1','1','1','1','0','1','0','0','0','1','1','0'),
            ('0','1','1','1','1','1','0','1','0','0','1','0','0','0'),
            ('0','1','1','1','1','1','0','1','0','0','1','0','1','0'),
            ('0','1','1','1','1','1','0','1','0','0','1','1','0','0'),
            ('0','1','1','1','1','1','0','1','0','0','1','1','1','0'),
            ('0','1','1','1','1','1','0','1','0','1','0','0','0','0'),
            ('0','1','1','1','1','1','0','1','0','1','0','0','1','0'),
            ('0','1','1','1','1','1','0','1','0','1','0','1','0','0'),
            ('0','1','1','1','1','1','0','1','0','1','0','1','1','0'),
            ('0','1','1','1','1','1','0','1','0','1','1','0','0','0'),
            ('0','1','1','1','1','1','0','1','0','1','1','0','1','0'),
            ('0','1','1','1','1','1','0','1','0','1','1','1','0','0'),
            ('0','1','1','1','1','1','0','1','0','1','1','1','1','0'),
            ('0','1','1','1','1','1','0','1','1','0','0','0','0','0'),
            ('0','1','1','1','1','1','0','1','1','0','0','0','1','0'),
            ('0','1','1','1','1','1','0','1','1','0','0','1','0','0'),
            ('0','1','1','1','1','1','0','1','1','0','0','1','1','0'),
            ('0','1','1','1','1','1','0','1','1','0','1','0','0','0'),
            ('0','1','1','1','1','1','0','1','1','0','1','0','1','0'),
            ('0','1','1','1','1','1','0','1','1','0','1','1','0','0'),
            ('0','1','1','1','1','1','0','1','1','0','1','1','1','0'),
            ('0','1','1','1','1','1','0','1','1','1','0','0','0','0'),
            ('0','1','1','1','1','1','0','1','1','1','0','0','1','0'),
            ('0','1','1','1','1','1','0','1','1','1','0','1','0','0'),
            ('0','1','1','1','1','1','0','1','1','1','0','1','1','0'),
            ('0','1','1','1','1','1','0','1','1','1','1','0','0','0'),
            ('0','1','1','1','1','1','0','1','1','1','1','0','1','0'),
            ('0','1','1','1','1','1','0','1','1','1','1','1','0','0'),
            ('0','1','1','1','1','1','0','1','1','1','1','1','1','0'),
            ('0','1','1','1','1','1','1','0','0','0','0','0','0','0'),
            ('0','1','1','1','1','1','1','0','0','0','0','0','1','0'),
            ('0','1','1','1','1','1','1','0','0','0','0','1','0','0'),
            ('0','1','1','1','1','1','1','0','0','0','0','1','1','0'),
            ('0','1','1','1','1','1','1','0','0','0','1','0','0','0'),
            ('0','1','1','1','1','1','1','0','0','0','1','0','1','0'),
            ('0','1','1','1','1','1','1','0','0','0','1','1','0','0'),
            ('0','1','1','1','1','1','1','0','0','0','1','1','1','0'),
            ('0','1','1','1','1','1','1','0','0','1','0','0','0','0'),
            ('0','1','1','1','1','1','1','0','0','1','0','0','1','0'),
            ('0','1','1','1','1','1','1','0','0','1','0','1','0','0'),
            ('0','1','1','1','1','1','1','0','0','1','0','1','1','0'),
            ('0','1','1','1','1','1','1','0','0','1','1','0','0','0'),
            ('0','1','1','1','1','1','1','0','0','1','1','0','1','0'),
            ('0','1','1','1','1','1','1','0','0','1','1','1','0','0'),
            ('0','1','1','1','1','1','1','0','0','1','1','1','1','0'),
            ('0','1','1','1','1','1','1','0','1','0','0','0','0','0'),
            ('0','1','1','1','1','1','1','0','1','0','0','0','1','0'),
            ('0','1','1','1','1','1','1','0','1','0','0','1','0','0'),
            ('0','1','1','1','1','1','1','0','1','0','0','1','1','0'),
            ('0','1','1','1','1','1','1','0','1','0','1','0','0','0'),
            ('0','1','1','1','1','1','1','0','1','0','1','0','1','0'),
            ('0','1','1','1','1','1','1','0','1','0','1','1','0','0'),
            ('0','1','1','1','1','1','1','0','1','0','1','1','1','0'),
            ('0','1','1','1','1','1','1','0','1','1','0','0','0','0'),
            ('0','1','1','1','1','1','1','0','1','1','0','0','1','0'),
            ('0','1','1','1','1','1','1','0','1','1','0','1','0','0'),
            ('0','1','1','1','1','1','1','0','1','1','0','1','1','0'),
            ('0','1','1','1','1','1','1','0','1','1','1','0','0','0'),
            ('0','1','1','1','1','1','1','0','1','1','1','0','1','0'),
            ('0','1','1','1','1','1','1','0','1','1','1','1','0','0'),
            ('0','1','1','1','1','1','1','0','1','1','1','1','1','0'),
            ('0','1','1','1','1','1','1','1','0','0','0','0','0','0'),
            ('0','1','1','1','1','1','1','1','0','0','0','0','1','0'),
            ('0','1','1','1','1','1','1','1','0','0','0','1','0','0'),
            ('0','1','1','1','1','1','1','1','0','0','0','1','1','0'),
            ('0','1','1','1','1','1','1','1','0','0','1','0','0','0'),
            ('0','1','1','1','1','1','1','1','0','0','1','0','1','0'),
            ('0','1','1','1','1','1','1','1','0','0','1','1','0','0'),
            ('0','1','1','1','1','1','1','1','0','0','1','1','1','0'),
            ('0','1','1','1','1','1','1','1','0','1','0','0','0','0'),
            ('0','1','1','1','1','1','1','1','0','1','0','0','1','0'),
            ('0','1','1','1','1','1','1','1','0','1','0','1','0','0'),
            ('0','1','1','1','1','1','1','1','0','1','0','1','1','0'),
            ('0','1','1','1','1','1','1','1','0','1','1','0','0','0'),
            ('0','1','1','1','1','1','1','1','0','1','1','0','1','0'),
            ('0','1','1','1','1','1','1','1','0','1','1','1','0','0'),
            ('0','1','1','1','1','1','1','1','0','1','1','1','1','0'),
            ('0','1','1','1','1','1','1','1','1','0','0','0','0','0'),
            ('0','1','1','1','1','1','1','1','1','0','0','0','1','0'),
            ('0','1','1','1','1','1','1','1','1','0','0','1','0','0'),
            ('0','1','1','1','1','1','1','1','1','0','0','1','1','0'),
            ('0','1','1','1','1','1','1','1','1','0','1','0','0','0'),
            ('0','1','1','1','1','1','1','1','1','0','1','0','1','0'),
            ('0','1','1','1','1','1','1','1','1','0','1','1','0','0'),
            ('0','1','1','1','1','1','1','1','1','0','1','1','1','0'),
            ('0','1','1','1','1','1','1','1','1','1','0','0','0','0'),
            ('0','1','1','1','1','1','1','1','1','1','0','0','1','0'),
            ('0','1','1','1','1','1','1','1','1','1','0','1','0','0'),
            ('0','1','1','1','1','1','1','1','1','1','0','1','1','0'),
            ('0','1','1','1','1','1','1','1','1','1','1','0','0','0'),
            ('0','1','1','1','1','1','1','1','1','1','1','0','1','0'),
            ('0','1','1','1','1','1','1','1','1','1','1','1','0','0'),
            ('0','1','1','1','1','1','1','1','1','1','1','1','1','0'),
            ('1','0','0','0','0','0','0','0','0','0','0','0','0','0'),
            ('1','0','0','0','0','0','0','0','0','0','0','0','1','0'),
            ('1','0','0','0','0','0','0','0','0','0','0','1','0','0'),
            ('1','0','0','0','0','0','0','0','0','0','0','1','1','0'),
            ('1','0','0','0','0','0','0','0','0','0','1','0','0','0'),
            ('1','0','0','0','0','0','0','0','0','0','1','0','1','0'),
            ('1','0','0','0','0','0','0','0','0','0','1','1','0','0'),
            ('1','0','0','0','0','0','0','0','0','0','1','1','1','0'),
            ('1','0','0','0','0','0','0','0','0','1','0','0','0','0'),
            ('1','0','0','0','0','0','0','0','0','1','0','0','1','0'),
            ('1','0','0','0','0','0','0','0','0','1','0','1','0','0'),
            ('1','0','0','0','0','0','0','0','0','1','0','1','1','0'),
            ('1','0','0','0','0','0','0','0','0','1','1','0','0','0'),
            ('1','0','0','0','0','0','0','0','0','1','1','0','1','0'),
            ('1','0','0','0','0','0','0','0','0','1','1','1','0','0'),
            ('1','0','0','0','0','0','0','0','0','1','1','1','1','0'),
            ('1','0','0','0','0','0','0','0','1','0','0','0','0','0'),
            ('1','0','0','0','0','0','0','0','1','0','0','0','1','0'),
            ('1','0','0','0','0','0','0','0','1','0','0','1','0','0'),
            ('1','0','0','0','0','0','0','0','1','0','0','1','1','0'),
            ('1','0','0','0','0','0','0','0','1','0','1','0','0','0'),
            ('1','0','0','0','0','0','0','0','1','0','1','0','1','0'),
            ('1','0','0','0','0','0','0','0','1','0','1','1','0','0'),
            ('1','0','0','0','0','0','0','0','1','0','1','1','1','0'),
            ('1','0','0','0','0','0','0','0','1','1','0','0','0','0'),
            ('1','0','0','0','0','0','0','0','1','1','0','0','1','0'),
            ('1','0','0','0','0','0','0','0','1','1','0','1','0','0'),
            ('1','0','0','0','0','0','0','0','1','1','0','1','1','0'),
            ('1','0','0','0','0','0','0','0','1','1','1','0','0','0'),
            ('1','0','0','0','0','0','0','0','1','1','1','0','1','0'),
            ('1','0','0','0','0','0','0','0','1','1','1','1','0','0'),
            ('1','0','0','0','0','0','0','0','1','1','1','1','1','0'),
            ('1','0','0','0','0','0','0','1','0','0','0','0','0','0'),
            ('1','0','0','0','0','0','0','1','0','0','0','0','1','0'),
            ('1','0','0','0','0','0','0','1','0','0','0','1','0','0'),
            ('1','0','0','0','0','0','0','1','0','0','0','1','1','0'),
            ('1','0','0','0','0','0','0','1','0','0','1','0','0','0'),
            ('1','0','0','0','0','0','0','1','0','0','1','0','1','0'),
            ('1','0','0','0','0','0','0','1','0','0','1','1','0','0'),
            ('1','0','0','0','0','0','0','1','0','0','1','1','1','0'),
            ('1','0','0','0','0','0','0','1','0','1','0','0','0','0'),
            ('1','0','0','0','0','0','0','1','0','1','0','0','1','0'),
            ('1','0','0','0','0','0','0','1','0','1','0','1','0','0'),
            ('1','0','0','0','0','0','0','1','0','1','0','1','1','0'),
            ('1','0','0','0','0','0','0','1','0','1','1','0','0','0'),
            ('1','0','0','0','0','0','0','1','0','1','1','0','1','0'),
            ('1','0','0','0','0','0','0','1','0','1','1','1','0','0'),
            ('1','0','0','0','0','0','0','1','0','1','1','1','1','0'),
            ('1','0','0','0','0','0','0','1','1','0','0','0','0','0'),
            ('1','0','0','0','0','0','0','1','1','0','0','0','1','0'),
            ('1','0','0','0','0','0','0','1','1','0','0','1','0','0'),
            ('1','0','0','0','0','0','0','1','1','0','0','1','1','0'),
            ('1','0','0','0','0','0','0','1','1','0','1','0','0','0'),
            ('1','0','0','0','0','0','0','1','1','0','1','0','1','0'),
            ('1','0','0','0','0','0','0','1','1','0','1','1','0','0'),
            ('1','0','0','0','0','0','0','1','1','0','1','1','1','0'),
            ('1','0','0','0','0','0','0','1','1','1','0','0','0','0'),
            ('1','0','0','0','0','0','0','1','1','1','0','0','1','0'),
            ('1','0','0','0','0','0','0','1','1','1','0','1','0','0'),
            ('1','0','0','0','0','0','0','1','1','1','0','1','1','0'),
            ('1','0','0','0','0','0','0','1','1','1','1','0','0','0'),
            ('1','0','0','0','0','0','0','1','1','1','1','0','1','0'),
            ('1','0','0','0','0','0','0','1','1','1','1','1','0','0'),
            ('1','0','0','0','0','0','0','1','1','1','1','1','1','0'),
            ('1','0','0','0','0','0','1','0','0','0','0','0','0','0'),
            ('1','0','0','0','0','0','1','0','0','0','0','0','1','0'),
            ('1','0','0','0','0','0','1','0','0','0','0','1','0','0'),
            ('1','0','0','0','0','0','1','0','0','0','0','1','1','0'),
            ('1','0','0','0','0','0','1','0','0','0','1','0','0','0'),
            ('1','0','0','0','0','0','1','0','0','0','1','0','1','0'),
            ('1','0','0','0','0','0','1','0','0','0','1','1','0','0'),
            ('1','0','0','0','0','0','1','0','0','0','1','1','1','0'),
            ('1','0','0','0','0','0','1','0','0','1','0','0','0','0'),
            ('1','0','0','0','0','0','1','0','0','1','0','0','1','0'),
            ('1','0','0','0','0','0','1','0','0','1','0','1','0','0'),
            ('1','0','0','0','0','0','1','0','0','1','0','1','1','0'),
            ('1','0','0','0','0','0','1','0','0','1','1','0','0','0'),
            ('1','0','0','0','0','0','1','0','0','1','1','0','1','0'),
            ('1','0','0','0','0','0','1','0','0','1','1','1','0','0'),
            ('1','0','0','0','0','0','1','0','0','1','1','1','1','0'),
            ('1','0','0','0','0','0','1','0','1','0','0','0','0','0'),
            ('1','0','0','0','0','0','1','0','1','0','0','0','1','0'),
            ('1','0','0','0','0','0','1','0','1','0','0','1','0','0'),
            ('1','0','0','0','0','0','1','0','1','0','0','1','1','0'),
            ('1','0','0','0','0','0','1','0','1','0','1','0','0','0'),
            ('1','0','0','0','0','0','1','0','1','0','1','0','1','0'),
            ('1','0','0','0','0','0','1','0','1','0','1','1','0','0'),
            ('1','0','0','0','0','0','1','0','1','0','1','1','1','0'),
            ('1','0','0','0','0','0','1','0','1','1','0','0','0','0'),
            ('1','0','0','0','0','0','1','0','1','1','0','0','1','0'),
            ('1','0','0','0','0','0','1','0','1','1','0','1','0','0'),
            ('1','0','0','0','0','0','1','0','1','1','0','1','1','0'),
            ('1','0','0','0','0','0','1','0','1','1','1','0','0','0'),
            ('1','0','0','0','0','0','1','0','1','1','1','0','1','0'),
            ('1','0','0','0','0','0','1','0','1','1','1','1','0','0'),
            ('1','0','0','0','0','0','1','0','1','1','1','1','1','0'),
            ('1','0','0','0','0','0','1','1','0','0','0','0','0','0'),
            ('1','0','0','0','0','0','1','1','0','0','0','0','1','0'),
            ('1','0','0','0','0','0','1','1','0','0','0','1','0','0'),
            ('1','0','0','0','0','0','1','1','0','0','0','1','1','0'),
            ('1','0','0','0','0','0','1','1','0','0','1','0','0','0'),
            ('1','0','0','0','0','0','1','1','0','0','1','0','1','0'),
            ('1','0','0','0','0','0','1','1','0','0','1','1','0','0'),
            ('1','0','0','0','0','0','1','1','0','0','1','1','1','0'),
            ('1','0','0','0','0','0','1','1','0','1','0','0','0','0'),
            ('1','0','0','0','0','0','1','1','0','1','0','0','1','0'),
            ('1','0','0','0','0','0','1','1','0','1','0','1','0','0'),
            ('1','0','0','0','0','0','1','1','0','1','0','1','1','0'),
            ('1','0','0','0','0','0','1','1','0','1','1','0','0','0'),
            ('1','0','0','0','0','0','1','1','0','1','1','0','1','0'),
            ('1','0','0','0','0','0','1','1','0','1','1','1','0','0'),
            ('1','0','0','0','0','0','1','1','0','1','1','1','1','0'),
            ('1','0','0','0','0','0','1','1','1','0','0','0','0','0'),
            ('1','0','0','0','0','0','1','1','1','0','0','0','1','0'),
            ('1','0','0','0','0','0','1','1','1','0','0','1','0','0'),
            ('1','0','0','0','0','0','1','1','1','0','0','1','1','0'),
            ('1','0','0','0','0','0','1','1','1','0','1','0','0','0'),
            ('1','0','0','0','0','0','1','1','1','0','1','0','1','0'),
            ('1','0','0','0','0','0','1','1','1','0','1','1','0','0'),
            ('1','0','0','0','0','0','1','1','1','0','1','1','1','0'),
            ('1','0','0','0','0','0','1','1','1','1','0','0','0','0'),
            ('1','0','0','0','0','0','1','1','1','1','0','0','1','0'),
            ('1','0','0','0','0','0','1','1','1','1','0','1','0','0'),
            ('1','0','0','0','0','0','1','1','1','1','0','1','1','0'),
            ('1','0','0','0','0','0','1','1','1','1','1','0','0','0'),
            ('1','0','0','0','0','0','1','1','1','1','1','0','1','0'),
            ('1','0','0','0','0','0','1','1','1','1','1','1','0','0'),
            ('1','0','0','0','0','0','1','1','1','1','1','1','1','0'),
            ('1','0','0','0','0','1','0','0','0','0','0','0','0','0'),
            ('1','0','0','0','0','1','0','0','0','0','0','0','1','0'),
            ('1','0','0','0','0','1','0','0','0','0','0','1','0','0'),
            ('1','0','0','0','0','1','0','0','0','0','0','1','1','0'),
            ('1','0','0','0','0','1','0','0','0','0','1','0','0','0'),
            ('1','0','0','0','0','1','0','0','0','0','1','0','1','0'),
            ('1','0','0','0','0','1','0','0','0','0','1','1','0','0'),
            ('1','0','0','0','0','1','0','0','0','0','1','1','1','0'),
            ('1','0','0','0','0','1','0','0','0','1','0','0','0','0'),
            ('1','0','0','0','0','1','0','0','0','1','0','0','1','0'),
            ('1','0','0','0','0','1','0','0','0','1','0','1','0','0'),
            ('1','0','0','0','0','1','0','0','0','1','0','1','1','0'),
            ('1','0','0','0','0','1','0','0','0','1','1','0','0','0'),
            ('1','0','0','0','0','1','0','0','0','1','1','0','1','0'),
            ('1','0','0','0','0','1','0','0','0','1','1','1','0','0'),
            ('1','0','0','0','0','1','0','0','0','1','1','1','1','0'),
            ('1','0','0','0','0','1','0','0','1','0','0','0','0','0'),
            ('1','0','0','0','0','1','0','0','1','0','0','0','1','0'),
            ('1','0','0','0','0','1','0','0','1','0','0','1','0','0'),
            ('1','0','0','0','0','1','0','0','1','0','0','1','1','0'),
            ('1','0','0','0','0','1','0','0','1','0','1','0','0','0'),
            ('1','0','0','0','0','1','0','0','1','0','1','0','1','0'),
            ('1','0','0','0','0','1','0','0','1','0','1','1','0','0'),
            ('1','0','0','0','0','1','0','0','1','0','1','1','1','0'),
            ('1','0','0','0','0','1','0','0','1','1','0','0','0','0'),
            ('1','0','0','0','0','1','0','0','1','1','0','0','1','0'),
            ('1','0','0','0','0','1','0','0','1','1','0','1','0','0'),
            ('1','0','0','0','0','1','0','0','1','1','0','1','1','0'),
            ('1','0','0','0','0','1','0','0','1','1','1','0','0','0'),
            ('1','0','0','0','0','1','0','0','1','1','1','0','1','0'),
            ('1','0','0','0','0','1','0','0','1','1','1','1','0','0'),
            ('1','0','0','0','0','1','0','0','1','1','1','1','1','0'),
            ('1','0','0','0','0','1','0','1','0','0','0','0','0','0'),
            ('1','0','0','0','0','1','0','1','0','0','0','0','1','0'),
            ('1','0','0','0','0','1','0','1','0','0','0','1','0','0'),
            ('1','0','0','0','0','1','0','1','0','0','0','1','1','0'),
            ('1','0','0','0','0','1','0','1','0','0','1','0','0','0'),
            ('1','0','0','0','0','1','0','1','0','0','1','0','1','0'),
            ('1','0','0','0','0','1','0','1','0','0','1','1','0','0'),
            ('1','0','0','0','0','1','0','1','0','0','1','1','1','0'),
            ('1','0','0','0','0','1','0','1','0','1','0','0','0','0'),
            ('1','0','0','0','0','1','0','1','0','1','0','0','1','0'),
            ('1','0','0','0','0','1','0','1','0','1','0','1','0','0'),
            ('1','0','0','0','0','1','0','1','0','1','0','1','1','0'),
            ('1','0','0','0','0','1','0','1','0','1','1','0','0','0'),
            ('1','0','0','0','0','1','0','1','0','1','1','0','1','0'),
            ('1','0','0','0','0','1','0','1','0','1','1','1','0','0'),
            ('1','0','0','0','0','1','0','1','0','1','1','1','1','0'),
            ('1','0','0','0','0','1','0','1','1','0','0','0','0','0'),
            ('1','0','0','0','0','1','0','1','1','0','0','0','1','0'),
            ('1','0','0','0','0','1','0','1','1','0','0','1','0','0'),
            ('1','0','0','0','0','1','0','1','1','0','0','1','1','0'),
            ('1','0','0','0','0','1','0','1','1','0','1','0','0','0'),
            ('1','0','0','0','0','1','0','1','1','0','1','0','1','0'),
            ('1','0','0','0','0','1','0','1','1','0','1','1','0','0'),
            ('1','0','0','0','0','1','0','1','1','0','1','1','1','0'),
            ('1','0','0','0','0','1','0','1','1','1','0','0','0','0'),
            ('1','0','0','0','0','1','0','1','1','1','0','0','1','0'),
            ('1','0','0','0','0','1','0','1','1','1','0','1','0','0'),
            ('1','0','0','0','0','1','0','1','1','1','0','1','1','0'),
            ('1','0','0','0','0','1','0','1','1','1','1','0','0','0'),
            ('1','0','0','0','0','1','0','1','1','1','1','0','1','0'),
            ('1','0','0','0','0','1','0','1','1','1','1','1','0','0'),
            ('1','0','0','0','0','1','0','1','1','1','1','1','1','0'),
            ('1','0','0','0','0','1','1','0','0','0','0','0','0','0'),
            ('1','0','0','0','0','1','1','0','0','0','0','0','1','0'),
            ('1','0','0','0','0','1','1','0','0','0','0','1','0','0'),
            ('1','0','0','0','0','1','1','0','0','0','0','1','1','0'),
            ('1','0','0','0','0','1','1','0','0','0','1','0','0','0'),
            ('1','0','0','0','0','1','1','0','0','0','1','0','1','0'),
            ('1','0','0','0','0','1','1','0','0','0','1','1','0','0'),
            ('1','0','0','0','0','1','1','0','0','0','1','1','1','0'),
            ('1','0','0','0','0','1','1','0','0','1','0','0','0','0'),
            ('1','0','0','0','0','1','1','0','0','1','0','0','1','0'),
            ('1','0','0','0','0','1','1','0','0','1','0','1','0','0'),
            ('1','0','0','0','0','1','1','0','0','1','0','1','1','0'),
            ('1','0','0','0','0','1','1','0','0','1','1','0','0','0'),
            ('1','0','0','0','0','1','1','0','0','1','1','0','1','0'),
            ('1','0','0','0','0','1','1','0','0','1','1','1','0','0'),
            ('1','0','0','0','0','1','1','0','0','1','1','1','1','0'),
            ('1','0','0','0','0','1','1','0','1','0','0','0','0','0'),
            ('1','0','0','0','0','1','1','0','1','0','0','0','1','0'),
            ('1','0','0','0','0','1','1','0','1','0','0','1','0','0'),
            ('1','0','0','0','0','1','1','0','1','0','0','1','1','0'),
            ('1','0','0','0','0','1','1','0','1','0','1','0','0','0'),
            ('1','0','0','0','0','1','1','0','1','0','1','0','1','0'),
            ('1','0','0','0','0','1','1','0','1','0','1','1','0','0'),
            ('1','0','0','0','0','1','1','0','1','0','1','1','1','0'),
            ('1','0','0','0','0','1','1','0','1','1','0','0','0','0'),
            ('1','0','0','0','0','1','1','0','1','1','0','0','1','0'),
            ('1','0','0','0','0','1','1','0','1','1','0','1','0','0'),
            ('1','0','0','0','0','1','1','0','1','1','0','1','1','0'),
            ('1','0','0','0','0','1','1','0','1','1','1','0','0','0'),
            ('1','0','0','0','0','1','1','0','1','1','1','0','1','0'),
            ('1','0','0','0','0','1','1','0','1','1','1','1','0','0'),
            ('1','0','0','0','0','1','1','0','1','1','1','1','1','0'),
            ('1','0','0','0','0','1','1','1','0','0','0','0','0','0'),
            ('1','0','0','0','0','1','1','1','0','0','0','0','1','0'),
            ('1','0','0','0','0','1','1','1','0','0','0','1','0','0'),
            ('1','0','0','0','0','1','1','1','0','0','0','1','1','0'),
            ('1','0','0','0','0','1','1','1','0','0','1','0','0','0'),
            ('1','0','0','0','0','1','1','1','0','0','1','0','1','0'),
            ('1','0','0','0','0','1','1','1','0','0','1','1','0','0'),
            ('1','0','0','0','0','1','1','1','0','0','1','1','1','0'),
            ('1','0','0','0','0','1','1','1','0','1','0','0','0','0'),
            ('1','0','0','0','0','1','1','1','0','1','0','0','1','0'),
            ('1','0','0','0','0','1','1','1','0','1','0','1','0','0'),
            ('1','0','0','0','0','1','1','1','0','1','0','1','1','0'),
            ('1','0','0','0','0','1','1','1','0','1','1','0','0','0'),
            ('1','0','0','0','0','1','1','1','0','1','1','0','1','0'),
            ('1','0','0','0','0','1','1','1','0','1','1','1','0','0'),
            ('1','0','0','0','0','1','1','1','0','1','1','1','1','0'),
            ('1','0','0','0','0','1','1','1','1','0','0','0','0','0'),
            ('1','0','0','0','0','1','1','1','1','0','0','0','1','0'),
            ('1','0','0','0','0','1','1','1','1','0','0','1','0','0'),
            ('1','0','0','0','0','1','1','1','1','0','0','1','1','0'),
            ('1','0','0','0','0','1','1','1','1','0','1','0','0','0'),
            ('1','0','0','0','0','1','1','1','1','0','1','0','1','0'),
            ('1','0','0','0','0','1','1','1','1','0','1','1','0','0'),
            ('1','0','0','0','0','1','1','1','1','0','1','1','1','0'),
            ('1','0','0','0','0','1','1','1','1','1','0','0','0','0'),
            ('1','0','0','0','0','1','1','1','1','1','0','0','1','0'),
            ('1','0','0','0','0','1','1','1','1','1','0','1','0','0'),
            ('1','0','0','0','0','1','1','1','1','1','0','1','1','0'),
            ('1','0','0','0','0','1','1','1','1','1','1','0','0','0'),
            ('1','0','0','0','0','1','1','1','1','1','1','0','1','0'),
            ('1','0','0','0','0','1','1','1','1','1','1','1','0','0'),
            ('1','0','0','0','0','1','1','1','1','1','1','1','1','0'),
            ('1','0','0','0','1','0','0','0','0','0','0','0','0','0'),
            ('1','0','0','0','1','0','0','0','0','0','0','0','1','0'),
            ('1','0','0','0','1','0','0','0','0','0','0','1','0','0'),
            ('1','0','0','0','1','0','0','0','0','0','0','1','1','0'),
            ('1','0','0','0','1','0','0','0','0','0','1','0','0','0'),
            ('1','0','0','0','1','0','0','0','0','0','1','0','1','0'),
            ('1','0','0','0','1','0','0','0','0','0','1','1','0','0'),
            ('1','0','0','0','1','0','0','0','0','0','1','1','1','0'),
            ('1','0','0','0','1','0','0','0','0','1','0','0','0','0'),
            ('1','0','0','0','1','0','0','0','0','1','0','0','1','0'),
            ('1','0','0','0','1','0','0','0','0','1','0','1','0','0'),
            ('1','0','0','0','1','0','0','0','0','1','0','1','1','0'),
            ('1','0','0','0','1','0','0','0','0','1','1','0','0','0'),
            ('1','0','0','0','1','0','0','0','0','1','1','0','1','0'),
            ('1','0','0','0','1','0','0','0','0','1','1','1','0','0'),
            ('1','0','0','0','1','0','0','0','0','1','1','1','1','0'),
            ('1','0','0','0','1','0','0','0','1','0','0','0','0','0'),
            ('1','0','0','0','1','0','0','0','1','0','0','0','1','0'),
            ('1','0','0','0','1','0','0','0','1','0','0','1','0','0'),
            ('1','0','0','0','1','0','0','0','1','0','0','1','1','0'),
            ('1','0','0','0','1','0','0','0','1','0','1','0','0','0'),
            ('1','0','0','0','1','0','0','0','1','0','1','0','1','0'),
            ('1','0','0','0','1','0','0','0','1','0','1','1','0','0'),
            ('1','0','0','0','1','0','0','0','1','0','1','1','1','0'),
            ('1','0','0','0','1','0','0','0','1','1','0','0','0','0'),
            ('1','0','0','0','1','0','0','0','1','1','0','0','1','0'),
            ('1','0','0','0','1','0','0','0','1','1','0','1','0','0'),
            ('1','0','0','0','1','0','0','0','1','1','0','1','1','0'),
            ('1','0','0','0','1','0','0','0','1','1','1','0','0','0'),
            ('1','0','0','0','1','0','0','0','1','1','1','0','1','0'),
            ('1','0','0','0','1','0','0','0','1','1','1','1','0','0'),
            ('1','0','0','0','1','0','0','0','1','1','1','1','1','0'),
            ('1','0','0','0','1','0','0','1','0','0','0','0','0','0'),
            ('1','0','0','0','1','0','0','1','0','0','0','0','1','0'),
            ('1','0','0','0','1','0','0','1','0','0','0','1','0','0'),
            ('1','0','0','0','1','0','0','1','0','0','0','1','1','0'),
            ('1','0','0','0','1','0','0','1','0','0','1','0','0','0'),
            ('1','0','0','0','1','0','0','1','0','0','1','0','1','0'),
            ('1','0','0','0','1','0','0','1','0','0','1','1','0','0'),
            ('1','0','0','0','1','0','0','1','0','0','1','1','1','0'),
            ('1','0','0','0','1','0','0','1','0','1','0','0','0','0'),
            ('1','0','0','0','1','0','0','1','0','1','0','0','1','0'),
            ('1','0','0','0','1','0','0','1','0','1','0','1','0','0'),
            ('1','0','0','0','1','0','0','1','0','1','0','1','1','0'),
            ('1','0','0','0','1','0','0','1','0','1','1','0','0','0'),
            ('1','0','0','0','1','0','0','1','0','1','1','0','1','0'),
            ('1','0','0','0','1','0','0','1','0','1','1','1','0','0'),
            ('1','0','0','0','1','0','0','1','0','1','1','1','1','0'),
            ('1','0','0','0','1','0','0','1','1','0','0','0','0','0'),
            ('1','0','0','0','1','0','0','1','1','0','0','0','1','0'),
            ('1','0','0','0','1','0','0','1','1','0','0','1','0','0'),
            ('1','0','0','0','1','0','0','1','1','0','0','1','1','0'),
            ('1','0','0','0','1','0','0','1','1','0','1','0','0','0'),
            ('1','0','0','0','1','0','0','1','1','0','1','0','1','0'),
            ('1','0','0','0','1','0','0','1','1','0','1','1','0','0'),
            ('1','0','0','0','1','0','0','1','1','0','1','1','1','0'),
            ('1','0','0','0','1','0','0','1','1','1','0','0','0','0'),
            ('1','0','0','0','1','0','0','1','1','1','0','0','1','0'),
            ('1','0','0','0','1','0','0','1','1','1','0','1','0','0'),
            ('1','0','0','0','1','0','0','1','1','1','0','1','1','0'),
            ('1','0','0','0','1','0','0','1','1','1','1','0','0','0'),
            ('1','0','0','0','1','0','0','1','1','1','1','0','1','0'),
            ('1','0','0','0','1','0','0','1','1','1','1','1','0','0'),
            ('1','0','0','0','1','0','0','1','1','1','1','1','1','0'),
            ('1','0','0','0','1','0','1','0','0','0','0','0','0','0'),
            ('1','0','0','0','1','0','1','0','0','0','0','0','1','0'),
            ('1','0','0','0','1','0','1','0','0','0','0','1','0','0'),
            ('1','0','0','0','1','0','1','0','0','0','0','1','1','0'),
            ('1','0','0','0','1','0','1','0','0','0','1','0','0','0'),
            ('1','0','0','0','1','0','1','0','0','0','1','0','1','0'),
            ('1','0','0','0','1','0','1','0','0','0','1','1','0','0'),
            ('1','0','0','0','1','0','1','0','0','0','1','1','1','0'),
            ('1','0','0','0','1','0','1','0','0','1','0','0','0','0'),
            ('1','0','0','0','1','0','1','0','0','1','0','0','1','0'),
            ('1','0','0','0','1','0','1','0','0','1','0','1','0','0'),
            ('1','0','0','0','1','0','1','0','0','1','0','1','1','0'),
            ('1','0','0','0','1','0','1','0','0','1','1','0','0','0'),
            ('1','0','0','0','1','0','1','0','0','1','1','0','1','0'),
            ('1','0','0','0','1','0','1','0','0','1','1','1','0','0'),
            ('1','0','0','0','1','0','1','0','0','1','1','1','1','0'),
            ('1','0','0','0','1','0','1','0','1','0','0','0','0','0'),
            ('1','0','0','0','1','0','1','0','1','0','0','0','1','0'),
            ('1','0','0','0','1','0','1','0','1','0','0','1','0','0'),
            ('1','0','0','0','1','0','1','0','1','0','0','1','1','0'),
            ('1','0','0','0','1','0','1','0','1','0','1','0','0','0'),
            ('1','0','0','0','1','0','1','0','1','0','1','0','1','0'),
            ('1','0','0','0','1','0','1','0','1','0','1','1','0','0'),
            ('1','0','0','0','1','0','1','0','1','0','1','1','1','0'),
            ('1','0','0','0','1','0','1','0','1','1','0','0','0','0'),
            ('1','0','0','0','1','0','1','0','1','1','0','0','1','0'),
            ('1','0','0','0','1','0','1','0','1','1','0','1','0','0'),
            ('1','0','0','0','1','0','1','0','1','1','0','1','1','0'),
            ('1','0','0','0','1','0','1','0','1','1','1','0','0','0'),
            ('1','0','0','0','1','0','1','0','1','1','1','0','1','0'),
            ('1','0','0','0','1','0','1','0','1','1','1','1','0','0'),
            ('1','0','0','0','1','0','1','0','1','1','1','1','1','0'),
            ('1','0','0','0','1','0','1','1','0','0','0','0','0','0'),
            ('1','0','0','0','1','0','1','1','0','0','0','0','1','0'),
            ('1','0','0','0','1','0','1','1','0','0','0','1','0','0'),
            ('1','0','0','0','1','0','1','1','0','0','0','1','1','0'),
            ('1','0','0','0','1','0','1','1','0','0','1','0','0','0'),
            ('1','0','0','0','1','0','1','1','0','0','1','0','1','0'),
            ('1','0','0','0','1','0','1','1','0','0','1','1','0','0'),
            ('1','0','0','0','1','0','1','1','0','0','1','1','1','0'),
            ('1','0','0','0','1','0','1','1','0','1','0','0','0','0'),
            ('1','0','0','0','1','0','1','1','0','1','0','0','1','0'),
            ('1','0','0','0','1','0','1','1','0','1','0','1','0','0'),
            ('1','0','0','0','1','0','1','1','0','1','0','1','1','0'),
            ('1','0','0','0','1','0','1','1','0','1','1','0','0','0'),
            ('1','0','0','0','1','0','1','1','0','1','1','0','1','0'),
            ('1','0','0','0','1','0','1','1','0','1','1','1','0','0'),
            ('1','0','0','0','1','0','1','1','0','1','1','1','1','0'),
            ('1','0','0','0','1','0','1','1','1','0','0','0','0','0'),
            ('1','0','0','0','1','0','1','1','1','0','0','0','1','0'),
            ('1','0','0','0','1','0','1','1','1','0','0','1','0','0'),
            ('1','0','0','0','1','0','1','1','1','0','0','1','1','0'),
            ('1','0','0','0','1','0','1','1','1','0','1','0','0','0'),
            ('1','0','0','0','1','0','1','1','1','0','1','0','1','0'),
            ('1','0','0','0','1','0','1','1','1','0','1','1','0','0'),
            ('1','0','0','0','1','0','1','1','1','0','1','1','1','0'),
            ('1','0','0','0','1','0','1','1','1','1','0','0','0','0'),
            ('1','0','0','0','1','0','1','1','1','1','0','0','1','0'),
            ('1','0','0','0','1','0','1','1','1','1','0','1','0','0'),
            ('1','0','0','0','1','0','1','1','1','1','0','1','1','0'),
            ('1','0','0','0','1','0','1','1','1','1','1','0','0','0'),
            ('1','0','0','0','1','0','1','1','1','1','1','0','1','0'),
            ('1','0','0','0','1','0','1','1','1','1','1','1','0','0'),
            ('1','0','0','0','1','0','1','1','1','1','1','1','1','0'),
            ('1','0','0','0','1','1','0','0','0','0','0','0','0','0'),
            ('1','0','0','0','1','1','0','0','0','0','0','0','1','0'),
            ('1','0','0','0','1','1','0','0','0','0','0','1','0','0'),
            ('1','0','0','0','1','1','0','0','0','0','0','1','1','0'),
            ('1','0','0','0','1','1','0','0','0','0','1','0','0','0'),
            ('1','0','0','0','1','1','0','0','0','0','1','0','1','0'),
            ('1','0','0','0','1','1','0','0','0','0','1','1','0','0'),
            ('1','0','0','0','1','1','0','0','0','0','1','1','1','0'),
            ('1','0','0','0','1','1','0','0','0','1','0','0','0','0'),
            ('1','0','0','0','1','1','0','0','0','1','0','0','1','0'),
            ('1','0','0','0','1','1','0','0','0','1','0','1','0','0'),
            ('1','0','0','0','1','1','0','0','0','1','0','1','1','0'),
            ('1','0','0','0','1','1','0','0','0','1','1','0','0','0'),
            ('1','0','0','0','1','1','0','0','0','1','1','0','1','0'),
            ('1','0','0','0','1','1','0','0','0','1','1','1','0','0'),
            ('1','0','0','0','1','1','0','0','0','1','1','1','1','0'),
            ('1','0','0','0','1','1','0','0','1','0','0','0','0','0'),
            ('1','0','0','0','1','1','0','0','1','0','0','0','1','0'),
            ('1','0','0','0','1','1','0','0','1','0','0','1','0','0'),
            ('1','0','0','0','1','1','0','0','1','0','0','1','1','0'),
            ('1','0','0','0','1','1','0','0','1','0','1','0','0','0'),
            ('1','0','0','0','1','1','0','0','1','0','1','0','1','0'),
            ('1','0','0','0','1','1','0','0','1','0','1','1','0','0'),
            ('1','0','0','0','1','1','0','0','1','0','1','1','1','0'),
            ('1','0','0','0','1','1','0','0','1','1','0','0','0','0'),
            ('1','0','0','0','1','1','0','0','1','1','0','0','1','0'),
            ('1','0','0','0','1','1','0','0','1','1','0','1','0','0'),
            ('1','0','0','0','1','1','0','0','1','1','0','1','1','0'),
            ('1','0','0','0','1','1','0','0','1','1','1','0','0','0'),
            ('1','0','0','0','1','1','0','0','1','1','1','0','1','0'),
            ('1','0','0','0','1','1','0','0','1','1','1','1','0','0'),
            ('1','0','0','0','1','1','0','0','1','1','1','1','1','0'),
            ('1','0','0','0','1','1','0','1','0','0','0','0','0','0'),
            ('1','0','0','0','1','1','0','1','0','0','0','0','1','0'),
            ('1','0','0','0','1','1','0','1','0','0','0','1','0','0'),
            ('1','0','0','0','1','1','0','1','0','0','0','1','1','0'),
            ('1','0','0','0','1','1','0','1','0','0','1','0','0','0'),
            ('1','0','0','0','1','1','0','1','0','0','1','0','1','0'),
            ('1','0','0','0','1','1','0','1','0','0','1','1','0','0'),
            ('1','0','0','0','1','1','0','1','0','0','1','1','1','0'),
            ('1','0','0','0','1','1','0','1','0','1','0','0','0','0'),
            ('1','0','0','0','1','1','0','1','0','1','0','0','1','0'),
            ('1','0','0','0','1','1','0','1','0','1','0','1','0','0'),
            ('1','0','0','0','1','1','0','1','0','1','0','1','1','0'),
            ('1','0','0','0','1','1','0','1','0','1','1','0','0','0'),
            ('1','0','0','0','1','1','0','1','0','1','1','0','1','0'),
            ('1','0','0','0','1','1','0','1','0','1','1','1','0','0'),
            ('1','0','0','0','1','1','0','1','0','1','1','1','1','0'),
            ('1','0','0','0','1','1','0','1','1','0','0','0','0','0'),
            ('1','0','0','0','1','1','0','1','1','0','0','0','1','0'),
            ('1','0','0','0','1','1','0','1','1','0','0','1','0','0'),
            ('1','0','0','0','1','1','0','1','1','0','0','1','1','0'),
            ('1','0','0','0','1','1','0','1','1','0','1','0','0','0'),
            ('1','0','0','0','1','1','0','1','1','0','1','0','1','0'),
            ('1','0','0','0','1','1','0','1','1','0','1','1','0','0'),
            ('1','0','0','0','1','1','0','1','1','0','1','1','1','0'),
            ('1','0','0','0','1','1','0','1','1','1','0','0','0','0'),
            ('1','0','0','0','1','1','0','1','1','1','0','0','1','0'),
            ('1','0','0','0','1','1','0','1','1','1','0','1','0','0'),
            ('1','0','0','0','1','1','0','1','1','1','0','1','1','0'),
            ('1','0','0','0','1','1','0','1','1','1','1','0','0','0'),
            ('1','0','0','0','1','1','0','1','1','1','1','0','1','0'),
            ('1','0','0','0','1','1','0','1','1','1','1','1','0','0'),
            ('1','0','0','0','1','1','0','1','1','1','1','1','1','0'),
            ('1','0','0','0','1','1','1','0','0','0','0','0','0','0'),
            ('1','0','0','0','1','1','1','0','0','0','0','0','1','0'),
            ('1','0','0','0','1','1','1','0','0','0','0','1','0','0'),
            ('1','0','0','0','1','1','1','0','0','0','0','1','1','0'),
            ('1','0','0','0','1','1','1','0','0','0','1','0','0','0'),
            ('1','0','0','0','1','1','1','0','0','0','1','0','1','0'),
            ('1','0','0','0','1','1','1','0','0','0','1','1','0','0'),
            ('1','0','0','0','1','1','1','0','0','0','1','1','1','0'),
            ('1','0','0','0','1','1','1','0','0','1','0','0','0','0'),
            ('1','0','0','0','1','1','1','0','0','1','0','0','1','0'),
            ('1','0','0','0','1','1','1','0','0','1','0','1','0','0'),
            ('1','0','0','0','1','1','1','0','0','1','0','1','1','0'),
            ('1','0','0','0','1','1','1','0','0','1','1','0','0','0'),
            ('1','0','0','0','1','1','1','0','0','1','1','0','1','0'),
            ('1','0','0','0','1','1','1','0','0','1','1','1','0','0'),
            ('1','0','0','0','1','1','1','0','0','1','1','1','1','0'),
            ('1','0','0','0','1','1','1','0','1','0','0','0','0','0'),
            ('1','0','0','0','1','1','1','0','1','0','0','0','1','0'),
            ('1','0','0','0','1','1','1','0','1','0','0','1','0','0'),
            ('1','0','0','0','1','1','1','0','1','0','0','1','1','0'),
            ('1','0','0','0','1','1','1','0','1','0','1','0','0','0'),
            ('1','0','0','0','1','1','1','0','1','0','1','0','1','0'),
            ('1','0','0','0','1','1','1','0','1','0','1','1','0','0'),
            ('1','0','0','0','1','1','1','0','1','0','1','1','1','0'),
            ('1','0','0','0','1','1','1','0','1','1','0','0','0','0'),
            ('1','0','0','0','1','1','1','0','1','1','0','0','1','0'),
            ('1','0','0','0','1','1','1','0','1','1','0','1','0','0'),
            ('1','0','0','0','1','1','1','0','1','1','0','1','1','0'),
            ('1','0','0','0','1','1','1','0','1','1','1','0','0','0'),
            ('1','0','0','0','1','1','1','0','1','1','1','0','1','0'),
            ('1','0','0','0','1','1','1','0','1','1','1','1','0','0'),
            ('1','0','0','0','1','1','1','0','1','1','1','1','1','0'),
            ('1','0','0','0','1','1','1','1','0','0','0','0','0','0'),
            ('1','0','0','0','1','1','1','1','0','0','0','0','1','0'),
            ('1','0','0','0','1','1','1','1','0','0','0','1','0','0'),
            ('1','0','0','0','1','1','1','1','0','0','0','1','1','0'),
            ('1','0','0','0','1','1','1','1','0','0','1','0','0','0'),
            ('1','0','0','0','1','1','1','1','0','0','1','0','1','0'),
            ('1','0','0','0','1','1','1','1','0','0','1','1','0','0'),
            ('1','0','0','0','1','1','1','1','0','0','1','1','1','0'),
            ('1','0','0','0','1','1','1','1','0','1','0','0','0','0'),
            ('1','0','0','0','1','1','1','1','0','1','0','0','1','0'),
            ('1','0','0','0','1','1','1','1','0','1','0','1','0','0'),
            ('1','0','0','0','1','1','1','1','0','1','0','1','1','0'),
            ('1','0','0','0','1','1','1','1','0','1','1','0','0','0'),
            ('1','0','0','0','1','1','1','1','0','1','1','0','1','0'),
            ('1','0','0','0','1','1','1','1','0','1','1','1','0','0'),
            ('1','0','0','0','1','1','1','1','0','1','1','1','1','0'),
            ('1','0','0','0','1','1','1','1','1','0','0','0','0','0'),
            ('1','0','0','0','1','1','1','1','1','0','0','0','1','0'),
            ('1','0','0','0','1','1','1','1','1','0','0','1','0','0'),
            ('1','0','0','0','1','1','1','1','1','0','0','1','1','0'),
            ('1','0','0','0','1','1','1','1','1','0','1','0','0','0'),
            ('1','0','0','0','1','1','1','1','1','0','1','0','1','0'),
            ('1','0','0','0','1','1','1','1','1','0','1','1','0','0'),
            ('1','0','0','0','1','1','1','1','1','0','1','1','1','0'),
            ('1','0','0','0','1','1','1','1','1','1','0','0','0','0'),
            ('1','0','0','0','1','1','1','1','1','1','0','0','1','0'),
            ('1','0','0','0','1','1','1','1','1','1','0','1','0','0'),
            ('1','0','0','0','1','1','1','1','1','1','0','1','1','0'),
            ('1','0','0','0','1','1','1','1','1','1','1','0','0','0'),
            ('1','0','0','0','1','1','1','1','1','1','1','0','1','0'),
            ('1','0','0','0','1','1','1','1','1','1','1','1','0','0'),
            ('1','0','0','0','1','1','1','1','1','1','1','1','1','0'),
            ('1','0','0','1','0','0','0','0','0','0','0','0','0','0'),
            ('1','0','0','1','0','0','0','0','0','0','0','0','1','0'),
            ('1','0','0','1','0','0','0','0','0','0','0','1','0','0'),
            ('1','0','0','1','0','0','0','0','0','0','0','1','1','0'),
            ('1','0','0','1','0','0','0','0','0','0','1','0','0','0'),
            ('1','0','0','1','0','0','0','0','0','0','1','0','1','0'),
            ('1','0','0','1','0','0','0','0','0','0','1','1','0','0'),
            ('1','0','0','1','0','0','0','0','0','0','1','1','1','0'),
            ('1','0','0','1','0','0','0','0','0','1','0','0','0','0'),
            ('1','0','0','1','0','0','0','0','0','1','0','0','1','0'),
            ('1','0','0','1','0','0','0','0','0','1','0','1','0','0'),
            ('1','0','0','1','0','0','0','0','0','1','0','1','1','0'),
            ('1','0','0','1','0','0','0','0','0','1','1','0','0','0'),
            ('1','0','0','1','0','0','0','0','0','1','1','0','1','0'),
            ('1','0','0','1','0','0','0','0','0','1','1','1','0','0'),
            ('1','0','0','1','0','0','0','0','0','1','1','1','1','0'),
            ('1','0','0','1','0','0','0','0','1','0','0','0','0','0'),
            ('1','0','0','1','0','0','0','0','1','0','0','0','1','0'),
            ('1','0','0','1','0','0','0','0','1','0','0','1','0','0'),
            ('1','0','0','1','0','0','0','0','1','0','0','1','1','0'),
            ('1','0','0','1','0','0','0','0','1','0','1','0','0','0'),
            ('1','0','0','1','0','0','0','0','1','0','1','0','1','0'),
            ('1','0','0','1','0','0','0','0','1','0','1','1','0','0'),
            ('1','0','0','1','0','0','0','0','1','0','1','1','1','0'),
            ('1','0','0','1','0','0','0','0','1','1','0','0','0','0'),
            ('1','0','0','1','0','0','0','0','1','1','0','0','1','0'),
            ('1','0','0','1','0','0','0','0','1','1','0','1','0','0'),
            ('1','0','0','1','0','0','0','0','1','1','0','1','1','0'),
            ('1','0','0','1','0','0','0','0','1','1','1','0','0','0'),
            ('1','0','0','1','0','0','0','0','1','1','1','0','1','0'),
            ('1','0','0','1','0','0','0','0','1','1','1','1','0','0'),
            ('1','0','0','1','0','0','0','0','1','1','1','1','1','0'),
            ('1','0','0','1','0','0','0','1','0','0','0','0','0','0'),
            ('1','0','0','1','0','0','0','1','0','0','0','0','1','0'),
            ('1','0','0','1','0','0','0','1','0','0','0','1','0','0'),
            ('1','0','0','1','0','0','0','1','0','0','0','1','1','0'),
            ('1','0','0','1','0','0','0','1','0','0','1','0','0','0'),
            ('1','0','0','1','0','0','0','1','0','0','1','0','1','0'),
            ('1','0','0','1','0','0','0','1','0','0','1','1','0','0'),
            ('1','0','0','1','0','0','0','1','0','0','1','1','1','0'),
            ('1','0','0','1','0','0','0','1','0','1','0','0','0','0'),
            ('1','0','0','1','0','0','0','1','0','1','0','0','1','0'),
            ('1','0','0','1','0','0','0','1','0','1','0','1','0','0'),
            ('1','0','0','1','0','0','0','1','0','1','0','1','1','0'),
            ('1','0','0','1','0','0','0','1','0','1','1','0','0','0'),
            ('1','0','0','1','0','0','0','1','0','1','1','0','1','0'),
            ('1','0','0','1','0','0','0','1','0','1','1','1','0','0'),
            ('1','0','0','1','0','0','0','1','0','1','1','1','1','0'),
            ('1','0','0','1','0','0','0','1','1','0','0','0','0','0'),
            ('1','0','0','1','0','0','0','1','1','0','0','0','1','0'),
            ('1','0','0','1','0','0','0','1','1','0','0','1','0','0'),
            ('1','0','0','1','0','0','0','1','1','0','0','1','1','0'),
            ('1','0','0','1','0','0','0','1','1','0','1','0','0','0'),
            ('1','0','0','1','0','0','0','1','1','0','1','0','1','0'),
            ('1','0','0','1','0','0','0','1','1','0','1','1','0','0'),
            ('1','0','0','1','0','0','0','1','1','0','1','1','1','0'),
            ('1','0','0','1','0','0','0','1','1','1','0','0','0','0'),
            ('1','0','0','1','0','0','0','1','1','1','0','0','1','0'),
            ('1','0','0','1','0','0','0','1','1','1','0','1','0','0'),
            ('1','0','0','1','0','0','0','1','1','1','0','1','1','0'),
            ('1','0','0','1','0','0','0','1','1','1','1','0','0','0'),
            ('1','0','0','1','0','0','0','1','1','1','1','0','1','0'),
            ('1','0','0','1','0','0','0','1','1','1','1','1','0','0'),
            ('1','0','0','1','0','0','0','1','1','1','1','1','1','0'),
            ('1','0','0','1','0','0','1','0','0','0','0','0','0','0'),
            ('1','0','0','1','0','0','1','0','0','0','0','0','1','0'),
            ('1','0','0','1','0','0','1','0','0','0','0','1','0','0'),
            ('1','0','0','1','0','0','1','0','0','0','0','1','1','0'),
            ('1','0','0','1','0','0','1','0','0','0','1','0','0','0'),
            ('1','0','0','1','0','0','1','0','0','0','1','0','1','0'),
            ('1','0','0','1','0','0','1','0','0','0','1','1','0','0'),
            ('1','0','0','1','0','0','1','0','0','0','1','1','1','0'),
            ('1','0','0','1','0','0','1','0','0','1','0','0','0','0'),
            ('1','0','0','1','0','0','1','0','0','1','0','0','1','0'),
            ('1','0','0','1','0','0','1','0','0','1','0','1','0','0'),
            ('1','0','0','1','0','0','1','0','0','1','0','1','1','0'),
            ('1','0','0','1','0','0','1','0','0','1','1','0','0','0'),
            ('1','0','0','1','0','0','1','0','0','1','1','0','1','0'),
            ('1','0','0','1','0','0','1','0','0','1','1','1','0','0'),
            ('1','0','0','1','0','0','1','0','0','1','1','1','1','0'),
            ('1','0','0','1','0','0','1','0','1','0','0','0','0','0'),
            ('1','0','0','1','0','0','1','0','1','0','0','0','1','0'),
            ('1','0','0','1','0','0','1','0','1','0','0','1','0','0'),
            ('1','0','0','1','0','0','1','0','1','0','0','1','1','0'),
            ('1','0','0','1','0','0','1','0','1','0','1','0','0','0'),
            ('1','0','0','1','0','0','1','0','1','0','1','0','1','0'),
            ('1','0','0','1','0','0','1','0','1','0','1','1','0','0'),
            ('1','0','0','1','0','0','1','0','1','0','1','1','1','0'),
            ('1','0','0','1','0','0','1','0','1','1','0','0','0','0'),
            ('1','0','0','1','0','0','1','0','1','1','0','0','1','0'),
            ('1','0','0','1','0','0','1','0','1','1','0','1','0','0'),
            ('1','0','0','1','0','0','1','0','1','1','0','1','1','0'),
            ('1','0','0','1','0','0','1','0','1','1','1','0','0','0'),
            ('1','0','0','1','0','0','1','0','1','1','1','0','1','0'),
            ('1','0','0','1','0','0','1','0','1','1','1','1','0','0'),
            ('1','0','0','1','0','0','1','0','1','1','1','1','1','0'),
            ('1','0','0','1','0','0','1','1','0','0','0','0','0','0'),
            ('1','0','0','1','0','0','1','1','0','0','0','0','1','0'),
            ('1','0','0','1','0','0','1','1','0','0','0','1','0','0'),
            ('1','0','0','1','0','0','1','1','0','0','0','1','1','0'),
            ('1','0','0','1','0','0','1','1','0','0','1','0','0','0'),
            ('1','0','0','1','0','0','1','1','0','0','1','0','1','0'),
            ('1','0','0','1','0','0','1','1','0','0','1','1','0','0'),
            ('1','0','0','1','0','0','1','1','0','0','1','1','1','0'),
            ('1','0','0','1','0','0','1','1','0','1','0','0','0','0'),
            ('1','0','0','1','0','0','1','1','0','1','0','0','1','0'),
            ('1','0','0','1','0','0','1','1','0','1','0','1','0','0'),
            ('1','0','0','1','0','0','1','1','0','1','0','1','1','0'),
            ('1','0','0','1','0','0','1','1','0','1','1','0','0','0'),
            ('1','0','0','1','0','0','1','1','0','1','1','0','1','0'),
            ('1','0','0','1','0','0','1','1','0','1','1','1','0','0'),
            ('1','0','0','1','0','0','1','1','0','1','1','1','1','0'),
            ('1','0','0','1','0','0','1','1','1','0','0','0','0','0'),
            ('1','0','0','1','0','0','1','1','1','0','0','0','1','0'),
            ('1','0','0','1','0','0','1','1','1','0','0','1','0','0'),
            ('1','0','0','1','0','0','1','1','1','0','0','1','1','0'),
            ('1','0','0','1','0','0','1','1','1','0','1','0','0','0'),
            ('1','0','0','1','0','0','1','1','1','0','1','0','1','0'),
            ('1','0','0','1','0','0','1','1','1','0','1','1','0','0'),
            ('1','0','0','1','0','0','1','1','1','0','1','1','1','0'),
            ('1','0','0','1','0','0','1','1','1','1','0','0','0','0'),
            ('1','0','0','1','0','0','1','1','1','1','0','0','1','0'),
            ('1','0','0','1','0','0','1','1','1','1','0','1','0','0'),
            ('1','0','0','1','0','0','1','1','1','1','0','1','1','0'),
            ('1','0','0','1','0','0','1','1','1','1','1','0','0','0'),
            ('1','0','0','1','0','0','1','1','1','1','1','0','1','0'),
            ('1','0','0','1','0','0','1','1','1','1','1','1','0','0'),
            ('1','0','0','1','0','0','1','1','1','1','1','1','1','0'),
            ('1','0','0','1','0','1','0','0','0','0','0','0','0','0'),
            ('1','0','0','1','0','1','0','0','0','0','0','0','1','0'),
            ('1','0','0','1','0','1','0','0','0','0','0','1','0','0'),
            ('1','0','0','1','0','1','0','0','0','0','0','1','1','0'),
            ('1','0','0','1','0','1','0','0','0','0','1','0','0','0'),
            ('1','0','0','1','0','1','0','0','0','0','1','0','1','0'),
            ('1','0','0','1','0','1','0','0','0','0','1','1','0','0'),
            ('1','0','0','1','0','1','0','0','0','0','1','1','1','0'),
            ('1','0','0','1','0','1','0','0','0','1','0','0','0','0'),
            ('1','0','0','1','0','1','0','0','0','1','0','0','1','0'),
            ('1','0','0','1','0','1','0','0','0','1','0','1','0','0'),
            ('1','0','0','1','0','1','0','0','0','1','0','1','1','0'),
            ('1','0','0','1','0','1','0','0','0','1','1','0','0','0'),
            ('1','0','0','1','0','1','0','0','0','1','1','0','1','0'),
            ('1','0','0','1','0','1','0','0','0','1','1','1','0','0'),
            ('1','0','0','1','0','1','0','0','0','1','1','1','1','0'),
            ('1','0','0','1','0','1','0','0','1','0','0','0','0','0'),
            ('1','0','0','1','0','1','0','0','1','0','0','0','1','0'),
            ('1','0','0','1','0','1','0','0','1','0','0','1','0','0'),
            ('1','0','0','1','0','1','0','0','1','0','0','1','1','0'),
            ('1','0','0','1','0','1','0','0','1','0','1','0','0','0'),
            ('1','0','0','1','0','1','0','0','1','0','1','0','1','0'),
            ('1','0','0','1','0','1','0','0','1','0','1','1','0','0'),
            ('1','0','0','1','0','1','0','0','1','0','1','1','1','0'),
            ('1','0','0','1','0','1','0','0','1','1','0','0','0','0'),
            ('1','0','0','1','0','1','0','0','1','1','0','0','1','0'),
            ('1','0','0','1','0','1','0','0','1','1','0','1','0','0'),
            ('1','0','0','1','0','1','0','0','1','1','0','1','1','0'),
            ('1','0','0','1','0','1','0','0','1','1','1','0','0','0'),
            ('1','0','0','1','0','1','0','0','1','1','1','0','1','0'),
            ('1','0','0','1','0','1','0','0','1','1','1','1','0','0'),
            ('1','0','0','1','0','1','0','0','1','1','1','1','1','0'),
            ('1','0','0','1','0','1','0','1','0','0','0','0','0','0'),
            ('1','0','0','1','0','1','0','1','0','0','0','0','1','0'),
            ('1','0','0','1','0','1','0','1','0','0','0','1','0','0'),
            ('1','0','0','1','0','1','0','1','0','0','0','1','1','0'),
            ('1','0','0','1','0','1','0','1','0','0','1','0','0','0'),
            ('1','0','0','1','0','1','0','1','0','0','1','0','1','0'),
            ('1','0','0','1','0','1','0','1','0','0','1','1','0','0'),
            ('1','0','0','1','0','1','0','1','0','0','1','1','1','0'),
            ('1','0','0','1','0','1','0','1','0','1','0','0','0','0'),
            ('1','0','0','1','0','1','0','1','0','1','0','0','1','0'),
            ('1','0','0','1','0','1','0','1','0','1','0','1','0','0'),
            ('1','0','0','1','0','1','0','1','0','1','0','1','1','0'),
            ('1','0','0','1','0','1','0','1','0','1','1','0','0','0'),
            ('1','0','0','1','0','1','0','1','0','1','1','0','1','0'),
            ('1','0','0','1','0','1','0','1','0','1','1','1','0','0'),
            ('1','0','0','1','0','1','0','1','0','1','1','1','1','0'),
            ('1','0','0','1','0','1','0','1','1','0','0','0','0','0'),
            ('1','0','0','1','0','1','0','1','1','0','0','0','1','0'),
            ('1','0','0','1','0','1','0','1','1','0','0','1','0','0'),
            ('1','0','0','1','0','1','0','1','1','0','0','1','1','0'),
            ('1','0','0','1','0','1','0','1','1','0','1','0','0','0'),
            ('1','0','0','1','0','1','0','1','1','0','1','0','1','0'),
            ('1','0','0','1','0','1','0','1','1','0','1','1','0','0'),
            ('1','0','0','1','0','1','0','1','1','0','1','1','1','0'),
            ('1','0','0','1','0','1','0','1','1','1','0','0','0','0'),
            ('1','0','0','1','0','1','0','1','1','1','0','0','1','0'),
            ('1','0','0','1','0','1','0','1','1','1','0','1','0','0'),
            ('1','0','0','1','0','1','0','1','1','1','0','1','1','0'),
            ('1','0','0','1','0','1','0','1','1','1','1','0','0','0'),
            ('1','0','0','1','0','1','0','1','1','1','1','0','1','0'),
            ('1','0','0','1','0','1','0','1','1','1','1','1','0','0'),
            ('1','0','0','1','0','1','0','1','1','1','1','1','1','0'),
            ('1','0','0','1','0','1','1','0','0','0','0','0','0','0'),
            ('1','0','0','1','0','1','1','0','0','0','0','0','1','0'),
            ('1','0','0','1','0','1','1','0','0','0','0','1','0','0'),
            ('1','0','0','1','0','1','1','0','0','0','0','1','1','0'),
            ('1','0','0','1','0','1','1','0','0','0','1','0','0','0'),
            ('1','0','0','1','0','1','1','0','0','0','1','0','1','0'),
            ('1','0','0','1','0','1','1','0','0','0','1','1','0','0'),
            ('1','0','0','1','0','1','1','0','0','0','1','1','1','0'),
            ('1','0','0','1','0','1','1','0','0','1','0','0','0','0'),
            ('1','0','0','1','0','1','1','0','0','1','0','0','1','0'),
            ('1','0','0','1','0','1','1','0','0','1','0','1','0','0'),
            ('1','0','0','1','0','1','1','0','0','1','0','1','1','0'),
            ('1','0','0','1','0','1','1','0','0','1','1','0','0','0'),
            ('1','0','0','1','0','1','1','0','0','1','1','0','1','0'),
            ('1','0','0','1','0','1','1','0','0','1','1','1','0','0'),
            ('1','0','0','1','0','1','1','0','0','1','1','1','1','0'),
            ('1','0','0','1','0','1','1','0','1','0','0','0','0','0'),
            ('1','0','0','1','0','1','1','0','1','0','0','0','1','0'),
            ('1','0','0','1','0','1','1','0','1','0','0','1','0','0'),
            ('1','0','0','1','0','1','1','0','1','0','0','1','1','0'),
            ('1','0','0','1','0','1','1','0','1','0','1','0','0','0'),
            ('1','0','0','1','0','1','1','0','1','0','1','0','1','0'),
            ('1','0','0','1','0','1','1','0','1','0','1','1','0','0'),
            ('1','0','0','1','0','1','1','0','1','0','1','1','1','0'),
            ('1','0','0','1','0','1','1','0','1','1','0','0','0','0'),
            ('1','0','0','1','0','1','1','0','1','1','0','0','1','0'),
            ('1','0','0','1','0','1','1','0','1','1','0','1','0','0'),
            ('1','0','0','1','0','1','1','0','1','1','0','1','1','0'),
            ('1','0','0','1','0','1','1','0','1','1','1','0','0','0'),
            ('1','0','0','1','0','1','1','0','1','1','1','0','1','0'),
            ('1','0','0','1','0','1','1','0','1','1','1','1','0','0'),
            ('1','0','0','1','0','1','1','0','1','1','1','1','1','0'),
            ('1','0','0','1','0','1','1','1','0','0','0','0','0','0'),
            ('1','0','0','1','0','1','1','1','0','0','0','0','1','0'),
            ('1','0','0','1','0','1','1','1','0','0','0','1','0','0'),
            ('1','0','0','1','0','1','1','1','0','0','0','1','1','0'),
            ('1','0','0','1','0','1','1','1','0','0','1','0','0','0'),
            ('1','0','0','1','0','1','1','1','0','0','1','0','1','0'),
            ('1','0','0','1','0','1','1','1','0','0','1','1','0','0'),
            ('1','0','0','1','0','1','1','1','0','0','1','1','1','0'),
            ('1','0','0','1','0','1','1','1','0','1','0','0','0','0'),
            ('1','0','0','1','0','1','1','1','0','1','0','0','1','0'),
            ('1','0','0','1','0','1','1','1','0','1','0','1','0','0'),
            ('1','0','0','1','0','1','1','1','0','1','0','1','1','0'),
            ('1','0','0','1','0','1','1','1','0','1','1','0','0','0'),
            ('1','0','0','1','0','1','1','1','0','1','1','0','1','0'),
            ('1','0','0','1','0','1','1','1','0','1','1','1','0','0'),
            ('1','0','0','1','0','1','1','1','0','1','1','1','1','0'),
            ('1','0','0','1','0','1','1','1','1','0','0','0','0','0'),
            ('1','0','0','1','0','1','1','1','1','0','0','0','1','0'),
            ('1','0','0','1','0','1','1','1','1','0','0','1','0','0'),
            ('1','0','0','1','0','1','1','1','1','0','0','1','1','0'),
            ('1','0','0','1','0','1','1','1','1','0','1','0','0','0'),
            ('1','0','0','1','0','1','1','1','1','0','1','0','1','0'),
            ('1','0','0','1','0','1','1','1','1','0','1','1','0','0'),
            ('1','0','0','1','0','1','1','1','1','0','1','1','1','0'),
            ('1','0','0','1','0','1','1','1','1','1','0','0','0','0'),
            ('1','0','0','1','0','1','1','1','1','1','0','0','1','0'),
            ('1','0','0','1','0','1','1','1','1','1','0','1','0','0'),
            ('1','0','0','1','0','1','1','1','1','1','0','1','1','0'),
            ('1','0','0','1','0','1','1','1','1','1','1','0','0','0'),
            ('1','0','0','1','0','1','1','1','1','1','1','0','1','0'),
            ('1','0','0','1','0','1','1','1','1','1','1','1','0','0'),
            ('1','0','0','1','0','1','1','1','1','1','1','1','1','0'),
            ('1','0','0','1','1','0','0','0','0','0','0','0','0','0'),
            ('1','0','0','1','1','0','0','0','0','0','0','0','1','0'),
            ('1','0','0','1','1','0','0','0','0','0','0','1','0','0'),
            ('1','0','0','1','1','0','0','0','0','0','0','1','1','0'),
            ('1','0','0','1','1','0','0','0','0','0','1','0','0','0'),
            ('1','0','0','1','1','0','0','0','0','0','1','0','1','0'),
            ('1','0','0','1','1','0','0','0','0','0','1','1','0','0'),
            ('1','0','0','1','1','0','0','0','0','0','1','1','1','0'),
            ('1','0','0','1','1','0','0','0','0','1','0','0','0','0'),
            ('1','0','0','1','1','0','0','0','0','1','0','0','1','0'),
            ('1','0','0','1','1','0','0','0','0','1','0','1','0','0'),
            ('1','0','0','1','1','0','0','0','0','1','0','1','1','0'),
            ('1','0','0','1','1','0','0','0','0','1','1','0','0','0'),
            ('1','0','0','1','1','0','0','0','0','1','1','0','1','0'),
            ('1','0','0','1','1','0','0','0','0','1','1','1','0','0'),
            ('1','0','0','1','1','0','0','0','0','1','1','1','1','0'),
            ('1','0','0','1','1','0','0','0','1','0','0','0','0','0'),
            ('1','0','0','1','1','0','0','0','1','0','0','0','1','0'),
            ('1','0','0','1','1','0','0','0','1','0','0','1','0','0'),
            ('1','0','0','1','1','0','0','0','1','0','0','1','1','0'),
            ('1','0','0','1','1','0','0','0','1','0','1','0','0','0'),
            ('1','0','0','1','1','0','0','0','1','0','1','0','1','0'),
            ('1','0','0','1','1','0','0','0','1','0','1','1','0','0'),
            ('1','0','0','1','1','0','0','0','1','0','1','1','1','0'),
            ('1','0','0','1','1','0','0','0','1','1','0','0','0','0'),
            ('1','0','0','1','1','0','0','0','1','1','0','0','1','0'),
            ('1','0','0','1','1','0','0','0','1','1','0','1','0','0'),
            ('1','0','0','1','1','0','0','0','1','1','0','1','1','0'),
            ('1','0','0','1','1','0','0','0','1','1','1','0','0','0'),
            ('1','0','0','1','1','0','0','0','1','1','1','0','1','0'),
            ('1','0','0','1','1','0','0','0','1','1','1','1','0','0'),
            ('1','0','0','1','1','0','0','0','1','1','1','1','1','0'),
            ('1','0','0','1','1','0','0','1','0','0','0','0','0','0'),
            ('1','0','0','1','1','0','0','1','0','0','0','0','1','0'),
            ('1','0','0','1','1','0','0','1','0','0','0','1','0','0'),
            ('1','0','0','1','1','0','0','1','0','0','0','1','1','0'),
            ('1','0','0','1','1','0','0','1','0','0','1','0','0','0'),
            ('1','0','0','1','1','0','0','1','0','0','1','0','1','0'),
            ('1','0','0','1','1','0','0','1','0','0','1','1','0','0'),
            ('1','0','0','1','1','0','0','1','0','0','1','1','1','0'),
            ('1','0','0','1','1','0','0','1','0','1','0','0','0','0'),
            ('1','0','0','1','1','0','0','1','0','1','0','0','1','0'),
            ('1','0','0','1','1','0','0','1','0','1','0','1','0','0'),
            ('1','0','0','1','1','0','0','1','0','1','0','1','1','0'),
            ('1','0','0','1','1','0','0','1','0','1','1','0','0','0'),
            ('1','0','0','1','1','0','0','1','0','1','1','0','1','0'),
            ('1','0','0','1','1','0','0','1','0','1','1','1','0','0'),
            ('1','0','0','1','1','0','0','1','0','1','1','1','1','0'),
            ('1','0','0','1','1','0','0','1','1','0','0','0','0','0'),
            ('1','0','0','1','1','0','0','1','1','0','0','0','1','0'),
            ('1','0','0','1','1','0','0','1','1','0','0','1','0','0'),
            ('1','0','0','1','1','0','0','1','1','0','0','1','1','0'),
            ('1','0','0','1','1','0','0','1','1','0','1','0','0','0'),
            ('1','0','0','1','1','0','0','1','1','0','1','0','1','0'),
            ('1','0','0','1','1','0','0','1','1','0','1','1','0','0'),
            ('1','0','0','1','1','0','0','1','1','0','1','1','1','0'),
            ('1','0','0','1','1','0','0','1','1','1','0','0','0','0'),
            ('1','0','0','1','1','0','0','1','1','1','0','0','1','0'),
            ('1','0','0','1','1','0','0','1','1','1','0','1','0','0'),
            ('1','0','0','1','1','0','0','1','1','1','0','1','1','0'),
            ('1','0','0','1','1','0','0','1','1','1','1','0','0','0'),
            ('1','0','0','1','1','0','0','1','1','1','1','0','1','0'),
            ('1','0','0','1','1','0','0','1','1','1','1','1','0','0'),
            ('1','0','0','1','1','0','0','1','1','1','1','1','1','0'),
            ('1','0','0','1','1','0','1','0','0','0','0','0','0','0'),
            ('1','0','0','1','1','0','1','0','0','0','0','0','1','0'),
            ('1','0','0','1','1','0','1','0','0','0','0','1','0','0'),
            ('1','0','0','1','1','0','1','0','0','0','0','1','1','0'),
            ('1','0','0','1','1','0','1','0','0','0','1','0','0','0'),
            ('1','0','0','1','1','0','1','0','0','0','1','0','1','0'),
            ('1','0','0','1','1','0','1','0','0','0','1','1','0','0'),
            ('1','0','0','1','1','0','1','0','0','0','1','1','1','0'),
            ('1','0','0','1','1','0','1','0','0','1','0','0','0','0'),
            ('1','0','0','1','1','0','1','0','0','1','0','0','1','0'),
            ('1','0','0','1','1','0','1','0','0','1','0','1','0','0'),
            ('1','0','0','1','1','0','1','0','0','1','0','1','1','0'),
            ('1','0','0','1','1','0','1','0','0','1','1','0','0','0'),
            ('1','0','0','1','1','0','1','0','0','1','1','0','1','0'),
            ('1','0','0','1','1','0','1','0','0','1','1','1','0','0'),
            ('1','0','0','1','1','0','1','0','0','1','1','1','1','0'),
            ('1','0','0','1','1','0','1','0','1','0','0','0','0','0'),
            ('1','0','0','1','1','0','1','0','1','0','0','0','1','0'),
            ('1','0','0','1','1','0','1','0','1','0','0','1','0','0'),
            ('1','0','0','1','1','0','1','0','1','0','0','1','1','0'),
            ('1','0','0','1','1','0','1','0','1','0','1','0','0','0'),
            ('1','0','0','1','1','0','1','0','1','0','1','0','1','0'),
            ('1','0','0','1','1','0','1','0','1','0','1','1','0','0'),
            ('1','0','0','1','1','0','1','0','1','0','1','1','1','0'),
            ('1','0','0','1','1','0','1','0','1','1','0','0','0','0'),
            ('1','0','0','1','1','0','1','0','1','1','0','0','1','0'),
            ('1','0','0','1','1','0','1','0','1','1','0','1','0','0'),
            ('1','0','0','1','1','0','1','0','1','1','0','1','1','0'),
            ('1','0','0','1','1','0','1','0','1','1','1','0','0','0'),
            ('1','0','0','1','1','0','1','0','1','1','1','0','1','0'),
            ('1','0','0','1','1','0','1','0','1','1','1','1','0','0'),
            ('1','0','0','1','1','0','1','0','1','1','1','1','1','0'),
            ('1','0','0','1','1','0','1','1','0','0','0','0','0','0'),
            ('1','0','0','1','1','0','1','1','0','0','0','0','1','0'),
            ('1','0','0','1','1','0','1','1','0','0','0','1','0','0'),
            ('1','0','0','1','1','0','1','1','0','0','0','1','1','0'),
            ('1','0','0','1','1','0','1','1','0','0','1','0','0','0'),
            ('1','0','0','1','1','0','1','1','0','0','1','0','1','0'),
            ('1','0','0','1','1','0','1','1','0','0','1','1','0','0'),
            ('1','0','0','1','1','0','1','1','0','0','1','1','1','0'),
            ('1','0','0','1','1','0','1','1','0','1','0','0','0','0'),
            ('1','0','0','1','1','0','1','1','0','1','0','0','1','0'),
            ('1','0','0','1','1','0','1','1','0','1','0','1','0','0'),
            ('1','0','0','1','1','0','1','1','0','1','0','1','1','0'),
            ('1','0','0','1','1','0','1','1','0','1','1','0','0','0'),
            ('1','0','0','1','1','0','1','1','0','1','1','0','1','0'),
            ('1','0','0','1','1','0','1','1','0','1','1','1','0','0'),
            ('1','0','0','1','1','0','1','1','0','1','1','1','1','0'),
            ('1','0','0','1','1','0','1','1','1','0','0','0','0','0'),
            ('1','0','0','1','1','0','1','1','1','0','0','0','1','0'),
            ('1','0','0','1','1','0','1','1','1','0','0','1','0','0'),
            ('1','0','0','1','1','0','1','1','1','0','0','1','1','0'),
            ('1','0','0','1','1','0','1','1','1','0','1','0','0','0'),
            ('1','0','0','1','1','0','1','1','1','0','1','0','1','0'),
            ('1','0','0','1','1','0','1','1','1','0','1','1','0','0'),
            ('1','0','0','1','1','0','1','1','1','0','1','1','1','0'),
            ('1','0','0','1','1','0','1','1','1','1','0','0','0','0'),
            ('1','0','0','1','1','0','1','1','1','1','0','0','1','0'),
            ('1','0','0','1','1','0','1','1','1','1','0','1','0','0'),
            ('1','0','0','1','1','0','1','1','1','1','0','1','1','0'),
            ('1','0','0','1','1','0','1','1','1','1','1','0','0','0'),
            ('1','0','0','1','1','0','1','1','1','1','1','0','1','0'),
            ('1','0','0','1','1','0','1','1','1','1','1','1','0','0'),
            ('1','0','0','1','1','0','1','1','1','1','1','1','1','0'),
            ('1','0','0','1','1','1','0','0','0','0','0','0','0','0'),
            ('1','0','0','1','1','1','0','0','0','0','0','0','1','0'),
            ('1','0','0','1','1','1','0','0','0','0','0','1','0','0'),
            ('1','0','0','1','1','1','0','0','0','0','0','1','1','0'),
            ('1','0','0','1','1','1','0','0','0','0','1','0','0','0'),
            ('1','0','0','1','1','1','0','0','0','0','1','0','1','0'),
            ('1','0','0','1','1','1','0','0','0','0','1','1','0','0'),
            ('1','0','0','1','1','1','0','0','0','0','1','1','1','0'),
            ('1','0','0','1','1','1','0','0','0','1','0','0','0','0'),
            ('1','0','0','1','1','1','0','0','0','1','0','0','1','0'),
            ('1','0','0','1','1','1','0','0','0','1','0','1','0','0'),
            ('1','0','0','1','1','1','0','0','0','1','0','1','1','0'),
            ('1','0','0','1','1','1','0','0','0','1','1','0','0','0'),
            ('1','0','0','1','1','1','0','0','0','1','1','0','1','0'),
            ('1','0','0','1','1','1','0','0','0','1','1','1','0','0'),
            ('1','0','0','1','1','1','0','0','0','1','1','1','1','0'),
            ('1','0','0','1','1','1','0','0','1','0','0','0','0','0'),
            ('1','0','0','1','1','1','0','0','1','0','0','0','1','0'),
            ('1','0','0','1','1','1','0','0','1','0','0','1','0','0'),
            ('1','0','0','1','1','1','0','0','1','0','0','1','1','0'),
            ('1','0','0','1','1','1','0','0','1','0','1','0','0','0'),
            ('1','0','0','1','1','1','0','0','1','0','1','0','1','0'),
            ('1','0','0','1','1','1','0','0','1','0','1','1','0','0'),
            ('1','0','0','1','1','1','0','0','1','0','1','1','1','0'),
            ('1','0','0','1','1','1','0','0','1','1','0','0','0','0'),
            ('1','0','0','1','1','1','0','0','1','1','0','0','1','0'),
            ('1','0','0','1','1','1','0','0','1','1','0','1','0','0'),
            ('1','0','0','1','1','1','0','0','1','1','0','1','1','0'),
            ('1','0','0','1','1','1','0','0','1','1','1','0','0','0'),
            ('1','0','0','1','1','1','0','0','1','1','1','0','1','0'),
            ('1','0','0','1','1','1','0','0','1','1','1','1','0','0'),
            ('1','0','0','1','1','1','0','0','1','1','1','1','1','0'),
            ('1','0','0','1','1','1','0','1','0','0','0','0','0','0'),
            ('1','0','0','1','1','1','0','1','0','0','0','0','1','0'),
            ('1','0','0','1','1','1','0','1','0','0','0','1','0','0'),
            ('1','0','0','1','1','1','0','1','0','0','0','1','1','0'),
            ('1','0','0','1','1','1','0','1','0','0','1','0','0','0'),
            ('1','0','0','1','1','1','0','1','0','0','1','0','1','0'),
            ('1','0','0','1','1','1','0','1','0','0','1','1','0','0'),
            ('1','0','0','1','1','1','0','1','0','0','1','1','1','0'),
            ('1','0','0','1','1','1','0','1','0','1','0','0','0','0'),
            ('1','0','0','1','1','1','0','1','0','1','0','0','1','0'),
            ('1','0','0','1','1','1','0','1','0','1','0','1','0','0'),
            ('1','0','0','1','1','1','0','1','0','1','0','1','1','0'),
            ('1','0','0','1','1','1','0','1','0','1','1','0','0','0'),
            ('1','0','0','1','1','1','0','1','0','1','1','0','1','0'),
            ('1','0','0','1','1','1','0','1','0','1','1','1','0','0'),
            ('1','0','0','1','1','1','0','1','0','1','1','1','1','0'),
            ('1','0','0','1','1','1','0','1','1','0','0','0','0','0'),
            ('1','0','0','1','1','1','0','1','1','0','0','0','1','0'),
            ('1','0','0','1','1','1','0','1','1','0','0','1','0','0'),
            ('1','0','0','1','1','1','0','1','1','0','0','1','1','0'),
            ('1','0','0','1','1','1','0','1','1','0','1','0','0','0'),
            ('1','0','0','1','1','1','0','1','1','0','1','0','1','0'),
            ('1','0','0','1','1','1','0','1','1','0','1','1','0','0'),
            ('1','0','0','1','1','1','0','1','1','0','1','1','1','0'),
            ('1','0','0','1','1','1','0','1','1','1','0','0','0','0'),
            ('1','0','0','1','1','1','0','1','1','1','0','0','1','0'),
            ('1','0','0','1','1','1','0','1','1','1','0','1','0','0'),
            ('1','0','0','1','1','1','0','1','1','1','0','1','1','0'),
            ('1','0','0','1','1','1','0','1','1','1','1','0','0','0'),
            ('1','0','0','1','1','1','0','1','1','1','1','0','1','0'),
            ('1','0','0','1','1','1','0','1','1','1','1','1','0','0'),
            ('1','0','0','1','1','1','0','1','1','1','1','1','1','0'),
            ('1','0','0','1','1','1','1','0','0','0','0','0','0','0'),
            ('1','0','0','1','1','1','1','0','0','0','0','0','1','0'),
            ('1','0','0','1','1','1','1','0','0','0','0','1','0','0'),
            ('1','0','0','1','1','1','1','0','0','0','0','1','1','0'),
            ('1','0','0','1','1','1','1','0','0','0','1','0','0','0'),
            ('1','0','0','1','1','1','1','0','0','0','1','0','1','0'),
            ('1','0','0','1','1','1','1','0','0','0','1','1','0','0'),
            ('1','0','0','1','1','1','1','0','0','0','1','1','1','0'),
            ('1','0','0','1','1','1','1','0','0','1','0','0','0','0'),
            ('1','0','0','1','1','1','1','0','0','1','0','0','1','0'),
            ('1','0','0','1','1','1','1','0','0','1','0','1','0','0'),
            ('1','0','0','1','1','1','1','0','0','1','0','1','1','0'),
            ('1','0','0','1','1','1','1','0','0','1','1','0','0','0'),
            ('1','0','0','1','1','1','1','0','0','1','1','0','1','0'),
            ('1','0','0','1','1','1','1','0','0','1','1','1','0','0'),
            ('1','0','0','1','1','1','1','0','0','1','1','1','1','0'),
            ('1','0','0','1','1','1','1','0','1','0','0','0','0','0'),
            ('1','0','0','1','1','1','1','0','1','0','0','0','1','0'),
            ('1','0','0','1','1','1','1','0','1','0','0','1','0','0'),
            ('1','0','0','1','1','1','1','0','1','0','0','1','1','0'),
            ('1','0','0','1','1','1','1','0','1','0','1','0','0','0'),
            ('1','0','0','1','1','1','1','0','1','0','1','0','1','0'),
            ('1','0','0','1','1','1','1','0','1','0','1','1','0','0'),
            ('1','0','0','1','1','1','1','0','1','0','1','1','1','0'),
            ('1','0','0','1','1','1','1','0','1','1','0','0','0','0'),
            ('1','0','0','1','1','1','1','0','1','1','0','0','1','0'),
            ('1','0','0','1','1','1','1','0','1','1','0','1','0','0'),
            ('1','0','0','1','1','1','1','0','1','1','0','1','1','0'),
            ('1','0','0','1','1','1','1','0','1','1','1','0','0','0'),
            ('1','0','0','1','1','1','1','0','1','1','1','0','1','0'),
            ('1','0','0','1','1','1','1','0','1','1','1','1','0','0'),
            ('1','0','0','1','1','1','1','0','1','1','1','1','1','0'),
            ('1','0','0','1','1','1','1','1','0','0','0','0','0','0'),
            ('1','0','0','1','1','1','1','1','0','0','0','0','1','0'),
            ('1','0','0','1','1','1','1','1','0','0','0','1','0','0'),
            ('1','0','0','1','1','1','1','1','0','0','0','1','1','0'),
            ('1','0','0','1','1','1','1','1','0','0','1','0','0','0'),
            ('1','0','0','1','1','1','1','1','0','0','1','0','1','0'),
            ('1','0','0','1','1','1','1','1','0','0','1','1','0','0'),
            ('1','0','0','1','1','1','1','1','0','0','1','1','1','0'),
            ('1','0','0','1','1','1','1','1','0','1','0','0','0','0'),
            ('1','0','0','1','1','1','1','1','0','1','0','0','1','0'),
            ('1','0','0','1','1','1','1','1','0','1','0','1','0','0'),
            ('1','0','0','1','1','1','1','1','0','1','0','1','1','0'),
            ('1','0','0','1','1','1','1','1','0','1','1','0','0','0'),
            ('1','0','0','1','1','1','1','1','0','1','1','0','1','0'),
            ('1','0','0','1','1','1','1','1','0','1','1','1','0','0'),
            ('1','0','0','1','1','1','1','1','0','1','1','1','1','0'),
            ('1','0','0','1','1','1','1','1','1','0','0','0','0','0'),
            ('1','0','0','1','1','1','1','1','1','0','0','0','1','0'),
            ('1','0','0','1','1','1','1','1','1','0','0','1','0','0'),
            ('1','0','0','1','1','1','1','1','1','0','0','1','1','0'),
            ('1','0','0','1','1','1','1','1','1','0','1','0','0','0'),
            ('1','0','0','1','1','1','1','1','1','0','1','0','1','0'),
            ('1','0','0','1','1','1','1','1','1','0','1','1','0','0'),
            ('1','0','0','1','1','1','1','1','1','0','1','1','1','0'),
            ('1','0','0','1','1','1','1','1','1','1','0','0','0','0'),
            ('1','0','0','1','1','1','1','1','1','1','0','0','1','0'),
            ('1','0','0','1','1','1','1','1','1','1','0','1','0','0'),
            ('1','0','0','1','1','1','1','1','1','1','0','1','1','0'),
            ('1','0','0','1','1','1','1','1','1','1','1','0','0','0'),
            ('1','0','0','1','1','1','1','1','1','1','1','0','1','0'),
            ('1','0','0','1','1','1','1','1','1','1','1','1','0','0'),
            ('1','0','0','1','1','1','1','1','1','1','1','1','1','0'),
            ('1','0','1','0','0','0','0','0','0','0','0','0','0','0'),
            ('1','0','1','0','0','0','0','0','0','0','0','0','1','0'),
            ('1','0','1','0','0','0','0','0','0','0','0','1','0','0'),
            ('1','0','1','0','0','0','0','0','0','0','0','1','1','0'),
            ('1','0','1','0','0','0','0','0','0','0','1','0','0','0'),
            ('1','0','1','0','0','0','0','0','0','0','1','0','1','0'),
            ('1','0','1','0','0','0','0','0','0','0','1','1','0','0'),
            ('1','0','1','0','0','0','0','0','0','0','1','1','1','0'),
            ('1','0','1','0','0','0','0','0','0','1','0','0','0','0'),
            ('1','0','1','0','0','0','0','0','0','1','0','0','1','0'),
            ('1','0','1','0','0','0','0','0','0','1','0','1','0','0'),
            ('1','0','1','0','0','0','0','0','0','1','0','1','1','0'),
            ('1','0','1','0','0','0','0','0','0','1','1','0','0','0'),
            ('1','0','1','0','0','0','0','0','0','1','1','0','1','0'),
            ('1','0','1','0','0','0','0','0','0','1','1','1','0','0'),
            ('1','0','1','0','0','0','0','0','0','1','1','1','1','0'),
            ('1','0','1','0','0','0','0','0','1','0','0','0','0','0'),
            ('1','0','1','0','0','0','0','0','1','0','0','0','1','0'),
            ('1','0','1','0','0','0','0','0','1','0','0','1','0','0'),
            ('1','0','1','0','0','0','0','0','1','0','0','1','1','0'),
            ('1','0','1','0','0','0','0','0','1','0','1','0','0','0'),
            ('1','0','1','0','0','0','0','0','1','0','1','0','1','0'),
            ('1','0','1','0','0','0','0','0','1','0','1','1','0','0'),
            ('1','0','1','0','0','0','0','0','1','0','1','1','1','0'),
            ('1','0','1','0','0','0','0','0','1','1','0','0','0','0'),
            ('1','0','1','0','0','0','0','0','1','1','0','0','1','0'),
            ('1','0','1','0','0','0','0','0','1','1','0','1','0','0'),
            ('1','0','1','0','0','0','0','0','1','1','0','1','1','0'),
            ('1','0','1','0','0','0','0','0','1','1','1','0','0','0'),
            ('1','0','1','0','0','0','0','0','1','1','1','0','1','0'),
            ('1','0','1','0','0','0','0','0','1','1','1','1','0','0'),
            ('1','0','1','0','0','0','0','0','1','1','1','1','1','0'),
            ('1','0','1','0','0','0','0','1','0','0','0','0','0','0'),
            ('1','0','1','0','0','0','0','1','0','0','0','0','1','0'),
            ('1','0','1','0','0','0','0','1','0','0','0','1','0','0'),
            ('1','0','1','0','0','0','0','1','0','0','0','1','1','0'),
            ('1','0','1','0','0','0','0','1','0','0','1','0','0','0'),
            ('1','0','1','0','0','0','0','1','0','0','1','0','1','0'),
            ('1','0','1','0','0','0','0','1','0','0','1','1','0','0'),
            ('1','0','1','0','0','0','0','1','0','0','1','1','1','0'),
            ('1','0','1','0','0','0','0','1','0','1','0','0','0','0'),
            ('1','0','1','0','0','0','0','1','0','1','0','0','1','0'),
            ('1','0','1','0','0','0','0','1','0','1','0','1','0','0'),
            ('1','0','1','0','0','0','0','1','0','1','0','1','1','0'),
            ('1','0','1','0','0','0','0','1','0','1','1','0','0','0'),
            ('1','0','1','0','0','0','0','1','0','1','1','0','1','0'),
            ('1','0','1','0','0','0','0','1','0','1','1','1','0','0'),
            ('1','0','1','0','0','0','0','1','0','1','1','1','1','0'),
            ('1','0','1','0','0','0','0','1','1','0','0','0','0','0'),
            ('1','0','1','0','0','0','0','1','1','0','0','0','1','0'),
            ('1','0','1','0','0','0','0','1','1','0','0','1','0','0'),
            ('1','0','1','0','0','0','0','1','1','0','0','1','1','0'),
            ('1','0','1','0','0','0','0','1','1','0','1','0','0','0'),
            ('1','0','1','0','0','0','0','1','1','0','1','0','1','0'),
            ('1','0','1','0','0','0','0','1','1','0','1','1','0','0'),
            ('1','0','1','0','0','0','0','1','1','0','1','1','1','0'),
            ('1','0','1','0','0','0','0','1','1','1','0','0','0','0'),
            ('1','0','1','0','0','0','0','1','1','1','0','0','1','0'),
            ('1','0','1','0','0','0','0','1','1','1','0','1','0','0'),
            ('1','0','1','0','0','0','0','1','1','1','0','1','1','0'),
            ('1','0','1','0','0','0','0','1','1','1','1','0','0','0'),
            ('1','0','1','0','0','0','0','1','1','1','1','0','1','0'),
            ('1','0','1','0','0','0','0','1','1','1','1','1','0','0'),
            ('1','0','1','0','0','0','0','1','1','1','1','1','1','0'),
            ('1','0','1','0','0','0','1','0','0','0','0','0','0','0'),
            ('1','0','1','0','0','0','1','0','0','0','0','0','1','0'),
            ('1','0','1','0','0','0','1','0','0','0','0','1','0','0'),
            ('1','0','1','0','0','0','1','0','0','0','0','1','1','0'),
            ('1','0','1','0','0','0','1','0','0','0','1','0','0','0'),
            ('1','0','1','0','0','0','1','0','0','0','1','0','1','0'),
            ('1','0','1','0','0','0','1','0','0','0','1','1','0','0'),
            ('1','0','1','0','0','0','1','0','0','0','1','1','1','0'),
            ('1','0','1','0','0','0','1','0','0','1','0','0','0','0'),
            ('1','0','1','0','0','0','1','0','0','1','0','0','1','0'),
            ('1','0','1','0','0','0','1','0','0','1','0','1','0','0'),
            ('1','0','1','0','0','0','1','0','0','1','0','1','1','0'),
            ('1','0','1','0','0','0','1','0','0','1','1','0','0','0'),
            ('1','0','1','0','0','0','1','0','0','1','1','0','1','0'),
            ('1','0','1','0','0','0','1','0','0','1','1','1','0','0'),
            ('1','0','1','0','0','0','1','0','0','1','1','1','1','0'),
            ('1','0','1','0','0','0','1','0','1','0','0','0','0','0'),
            ('1','0','1','0','0','0','1','0','1','0','0','0','1','0'),
            ('1','0','1','0','0','0','1','0','1','0','0','1','0','0'),
            ('1','0','1','0','0','0','1','0','1','0','0','1','1','0'),
            ('1','0','1','0','0','0','1','0','1','0','1','0','0','0'),
            ('1','0','1','0','0','0','1','0','1','0','1','0','1','0'),
            ('1','0','1','0','0','0','1','0','1','0','1','1','0','0'),
            ('1','0','1','0','0','0','1','0','1','0','1','1','1','0'),
            ('1','0','1','0','0','0','1','0','1','1','0','0','0','0'),
            ('1','0','1','0','0','0','1','0','1','1','0','0','1','0'),
            ('1','0','1','0','0','0','1','0','1','1','0','1','0','0'),
            ('1','0','1','0','0','0','1','0','1','1','0','1','1','0'),
            ('1','0','1','0','0','0','1','0','1','1','1','0','0','0'),
            ('1','0','1','0','0','0','1','0','1','1','1','0','1','0'),
            ('1','0','1','0','0','0','1','0','1','1','1','1','0','0'),
            ('1','0','1','0','0','0','1','0','1','1','1','1','1','0'),
            ('1','0','1','0','0','0','1','1','0','0','0','0','0','0'),
            ('1','0','1','0','0','0','1','1','0','0','0','0','1','0'),
            ('1','0','1','0','0','0','1','1','0','0','0','1','0','0'),
            ('1','0','1','0','0','0','1','1','0','0','0','1','1','0'),
            ('1','0','1','0','0','0','1','1','0','0','1','0','0','0'),
            ('1','0','1','0','0','0','1','1','0','0','1','0','1','0'),
            ('1','0','1','0','0','0','1','1','0','0','1','1','0','0'),
            ('1','0','1','0','0','0','1','1','0','0','1','1','1','0'),
            ('1','0','1','0','0','0','1','1','0','1','0','0','0','0'),
            ('1','0','1','0','0','0','1','1','0','1','0','0','1','0'),
            ('1','0','1','0','0','0','1','1','0','1','0','1','0','0'),
            ('1','0','1','0','0','0','1','1','0','1','0','1','1','0'),
            ('1','0','1','0','0','0','1','1','0','1','1','0','0','0'),
            ('1','0','1','0','0','0','1','1','0','1','1','0','1','0'),
            ('1','0','1','0','0','0','1','1','0','1','1','1','0','0'),
            ('1','0','1','0','0','0','1','1','0','1','1','1','1','0'),
            ('1','0','1','0','0','0','1','1','1','0','0','0','0','0'),
            ('1','0','1','0','0','0','1','1','1','0','0','0','1','0'),
            ('1','0','1','0','0','0','1','1','1','0','0','1','0','0'),
            ('1','0','1','0','0','0','1','1','1','0','0','1','1','0'),
            ('1','0','1','0','0','0','1','1','1','0','1','0','0','0'),
            ('1','0','1','0','0','0','1','1','1','0','1','0','1','0'),
            ('1','0','1','0','0','0','1','1','1','0','1','1','0','0'),
            ('1','0','1','0','0','0','1','1','1','0','1','1','1','0'),
            ('1','0','1','0','0','0','1','1','1','1','0','0','0','0'),
            ('1','0','1','0','0','0','1','1','1','1','0','0','1','0'),
            ('1','0','1','0','0','0','1','1','1','1','0','1','0','0'),
            ('1','0','1','0','0','0','1','1','1','1','0','1','1','0'),
            ('1','0','1','0','0','0','1','1','1','1','1','0','0','0'),
            ('1','0','1','0','0','0','1','1','1','1','1','0','1','0'),
            ('1','0','1','0','0','0','1','1','1','1','1','1','0','0'),
            ('1','0','1','0','0','0','1','1','1','1','1','1','1','0'),
            ('1','0','1','0','0','1','0','0','0','0','0','0','0','0'),
            ('1','0','1','0','0','1','0','0','0','0','0','0','1','0'),
            ('1','0','1','0','0','1','0','0','0','0','0','1','0','0'),
            ('1','0','1','0','0','1','0','0','0','0','0','1','1','0'),
            ('1','0','1','0','0','1','0','0','0','0','1','0','0','0'),
            ('1','0','1','0','0','1','0','0','0','0','1','0','1','0'),
            ('1','0','1','0','0','1','0','0','0','0','1','1','0','0'),
            ('1','0','1','0','0','1','0','0','0','0','1','1','1','0'),
            ('1','0','1','0','0','1','0','0','0','1','0','0','0','0'),
            ('1','0','1','0','0','1','0','0','0','1','0','0','1','0'),
            ('1','0','1','0','0','1','0','0','0','1','0','1','0','0'),
            ('1','0','1','0','0','1','0','0','0','1','0','1','1','0'),
            ('1','0','1','0','0','1','0','0','0','1','1','0','0','0'),
            ('1','0','1','0','0','1','0','0','0','1','1','0','1','0'),
            ('1','0','1','0','0','1','0','0','0','1','1','1','0','0'),
            ('1','0','1','0','0','1','0','0','0','1','1','1','1','0'),
            ('1','0','1','0','0','1','0','0','1','0','0','0','0','0'),
            ('1','0','1','0','0','1','0','0','1','0','0','0','1','0'),
            ('1','0','1','0','0','1','0','0','1','0','0','1','0','0'),
            ('1','0','1','0','0','1','0','0','1','0','0','1','1','0'),
            ('1','0','1','0','0','1','0','0','1','0','1','0','0','0'),
            ('1','0','1','0','0','1','0','0','1','0','1','0','1','0'),
            ('1','0','1','0','0','1','0','0','1','0','1','1','0','0'),
            ('1','0','1','0','0','1','0','0','1','0','1','1','1','0'),
            ('1','0','1','0','0','1','0','0','1','1','0','0','0','0'),
            ('1','0','1','0','0','1','0','0','1','1','0','0','1','0'),
            ('1','0','1','0','0','1','0','0','1','1','0','1','0','0'),
            ('1','0','1','0','0','1','0','0','1','1','0','1','1','0'),
            ('1','0','1','0','0','1','0','0','1','1','1','0','0','0'),
            ('1','0','1','0','0','1','0','0','1','1','1','0','1','0'),
            ('1','0','1','0','0','1','0','0','1','1','1','1','0','0'),
            ('1','0','1','0','0','1','0','0','1','1','1','1','1','0'),
            ('1','0','1','0','0','1','0','1','0','0','0','0','0','0'),
            ('1','0','1','0','0','1','0','1','0','0','0','0','1','0'),
            ('1','0','1','0','0','1','0','1','0','0','0','1','0','0'),
            ('1','0','1','0','0','1','0','1','0','0','0','1','1','0'),
            ('1','0','1','0','0','1','0','1','0','0','1','0','0','0'),
            ('1','0','1','0','0','1','0','1','0','0','1','0','1','0'),
            ('1','0','1','0','0','1','0','1','0','0','1','1','0','0'),
            ('1','0','1','0','0','1','0','1','0','0','1','1','1','0'),
            ('1','0','1','0','0','1','0','1','0','1','0','0','0','0'),
            ('1','0','1','0','0','1','0','1','0','1','0','0','1','0'),
            ('1','0','1','0','0','1','0','1','0','1','0','1','0','0'),
            ('1','0','1','0','0','1','0','1','0','1','0','1','1','0'),
            ('1','0','1','0','0','1','0','1','0','1','1','0','0','0'),
            ('1','0','1','0','0','1','0','1','0','1','1','0','1','0'),
            ('1','0','1','0','0','1','0','1','0','1','1','1','0','0'),
            ('1','0','1','0','0','1','0','1','0','1','1','1','1','0'),
            ('1','0','1','0','0','1','0','1','1','0','0','0','0','0'),
            ('1','0','1','0','0','1','0','1','1','0','0','0','1','0'),
            ('1','0','1','0','0','1','0','1','1','0','0','1','0','0'),
            ('1','0','1','0','0','1','0','1','1','0','0','1','1','0'),
            ('1','0','1','0','0','1','0','1','1','0','1','0','0','0'),
            ('1','0','1','0','0','1','0','1','1','0','1','0','1','0'),
            ('1','0','1','0','0','1','0','1','1','0','1','1','0','0'),
            ('1','0','1','0','0','1','0','1','1','0','1','1','1','0'),
            ('1','0','1','0','0','1','0','1','1','1','0','0','0','0'),
            ('1','0','1','0','0','1','0','1','1','1','0','0','1','0'),
            ('1','0','1','0','0','1','0','1','1','1','0','1','0','0'),
            ('1','0','1','0','0','1','0','1','1','1','0','1','1','0'),
            ('1','0','1','0','0','1','0','1','1','1','1','0','0','0'),
            ('1','0','1','0','0','1','0','1','1','1','1','0','1','0'),
            ('1','0','1','0','0','1','0','1','1','1','1','1','0','0'),
            ('1','0','1','0','0','1','0','1','1','1','1','1','1','0'),
            ('1','0','1','0','0','1','1','0','0','0','0','0','0','0'),
            ('1','0','1','0','0','1','1','0','0','0','0','0','1','0'),
            ('1','0','1','0','0','1','1','0','0','0','0','1','0','0'),
            ('1','0','1','0','0','1','1','0','0','0','0','1','1','0'),
            ('1','0','1','0','0','1','1','0','0','0','1','0','0','0'),
            ('1','0','1','0','0','1','1','0','0','0','1','0','1','0'),
            ('1','0','1','0','0','1','1','0','0','0','1','1','0','0'),
            ('1','0','1','0','0','1','1','0','0','0','1','1','1','0'),
            ('1','0','1','0','0','1','1','0','0','1','0','0','0','0'),
            ('1','0','1','0','0','1','1','0','0','1','0','0','1','0'),
            ('1','0','1','0','0','1','1','0','0','1','0','1','0','0'),
            ('1','0','1','0','0','1','1','0','0','1','0','1','1','0'),
            ('1','0','1','0','0','1','1','0','0','1','1','0','0','0'),
            ('1','0','1','0','0','1','1','0','0','1','1','0','1','0'),
            ('1','0','1','0','0','1','1','0','0','1','1','1','0','0'),
            ('1','0','1','0','0','1','1','0','0','1','1','1','1','0'),
            ('1','0','1','0','0','1','1','0','1','0','0','0','0','0'),
            ('1','0','1','0','0','1','1','0','1','0','0','0','1','0'),
            ('1','0','1','0','0','1','1','0','1','0','0','1','0','0'),
            ('1','0','1','0','0','1','1','0','1','0','0','1','1','0'),
            ('1','0','1','0','0','1','1','0','1','0','1','0','0','0'),
            ('1','0','1','0','0','1','1','0','1','0','1','0','1','0'),
            ('1','0','1','0','0','1','1','0','1','0','1','1','0','0'),
            ('1','0','1','0','0','1','1','0','1','0','1','1','1','0'),
            ('1','0','1','0','0','1','1','0','1','1','0','0','0','0'),
            ('1','0','1','0','0','1','1','0','1','1','0','0','1','0'),
            ('1','0','1','0','0','1','1','0','1','1','0','1','0','0'),
            ('1','0','1','0','0','1','1','0','1','1','0','1','1','0'),
            ('1','0','1','0','0','1','1','0','1','1','1','0','0','0'),
            ('1','0','1','0','0','1','1','0','1','1','1','0','1','0'),
            ('1','0','1','0','0','1','1','0','1','1','1','1','0','0'),
            ('1','0','1','0','0','1','1','0','1','1','1','1','1','0'),
            ('1','0','1','0','0','1','1','1','0','0','0','0','0','0'),
            ('1','0','1','0','0','1','1','1','0','0','0','0','1','0'),
            ('1','0','1','0','0','1','1','1','0','0','0','1','0','0'),
            ('1','0','1','0','0','1','1','1','0','0','0','1','1','0'),
            ('1','0','1','0','0','1','1','1','0','0','1','0','0','0'),
            ('1','0','1','0','0','1','1','1','0','0','1','0','1','0'),
            ('1','0','1','0','0','1','1','1','0','0','1','1','0','0'),
            ('1','0','1','0','0','1','1','1','0','0','1','1','1','0'),
            ('1','0','1','0','0','1','1','1','0','1','0','0','0','0'),
            ('1','0','1','0','0','1','1','1','0','1','0','0','1','0'),
            ('1','0','1','0','0','1','1','1','0','1','0','1','0','0'),
            ('1','0','1','0','0','1','1','1','0','1','0','1','1','0'),
            ('1','0','1','0','0','1','1','1','0','1','1','0','0','0'),
            ('1','0','1','0','0','1','1','1','0','1','1','0','1','0'),
            ('1','0','1','0','0','1','1','1','0','1','1','1','0','0'),
            ('1','0','1','0','0','1','1','1','0','1','1','1','1','0'),
            ('1','0','1','0','0','1','1','1','1','0','0','0','0','0'),
            ('1','0','1','0','0','1','1','1','1','0','0','0','1','0'),
            ('1','0','1','0','0','1','1','1','1','0','0','1','0','0'),
            ('1','0','1','0','0','1','1','1','1','0','0','1','1','0'),
            ('1','0','1','0','0','1','1','1','1','0','1','0','0','0'),
            ('1','0','1','0','0','1','1','1','1','0','1','0','1','0'),
            ('1','0','1','0','0','1','1','1','1','0','1','1','0','0'),
            ('1','0','1','0','0','1','1','1','1','0','1','1','1','0'),
            ('1','0','1','0','0','1','1','1','1','1','0','0','0','0'),
            ('1','0','1','0','0','1','1','1','1','1','0','0','1','0'),
            ('1','0','1','0','0','1','1','1','1','1','0','1','0','0'),
            ('1','0','1','0','0','1','1','1','1','1','0','1','1','0'),
            ('1','0','1','0','0','1','1','1','1','1','1','0','0','0'),
            ('1','0','1','0','0','1','1','1','1','1','1','0','1','0'),
            ('1','0','1','0','0','1','1','1','1','1','1','1','0','0'),
            ('1','0','1','0','0','1','1','1','1','1','1','1','1','0'),
            ('1','0','1','0','1','0','0','0','0','0','0','0','0','0'),
            ('1','0','1','0','1','0','0','0','0','0','0','0','1','0'),
            ('1','0','1','0','1','0','0','0','0','0','0','1','0','0'),
            ('1','0','1','0','1','0','0','0','0','0','0','1','1','0'),
            ('1','0','1','0','1','0','0','0','0','0','1','0','0','0'),
            ('1','0','1','0','1','0','0','0','0','0','1','0','1','0'),
            ('1','0','1','0','1','0','0','0','0','0','1','1','0','0'),
            ('1','0','1','0','1','0','0','0','0','0','1','1','1','0'),
            ('1','0','1','0','1','0','0','0','0','1','0','0','0','0'),
            ('1','0','1','0','1','0','0','0','0','1','0','0','1','0'),
            ('1','0','1','0','1','0','0','0','0','1','0','1','0','0'),
            ('1','0','1','0','1','0','0','0','0','1','0','1','1','0'),
            ('1','0','1','0','1','0','0','0','0','1','1','0','0','0'),
            ('1','0','1','0','1','0','0','0','0','1','1','0','1','0'),
            ('1','0','1','0','1','0','0','0','0','1','1','1','0','0'),
            ('1','0','1','0','1','0','0','0','0','1','1','1','1','0'),
            ('1','0','1','0','1','0','0','0','1','0','0','0','0','0'),
            ('1','0','1','0','1','0','0','0','1','0','0','0','1','0'),
            ('1','0','1','0','1','0','0','0','1','0','0','1','0','0'),
            ('1','0','1','0','1','0','0','0','1','0','0','1','1','0'),
            ('1','0','1','0','1','0','0','0','1','0','1','0','0','0'),
            ('1','0','1','0','1','0','0','0','1','0','1','0','1','0'),
            ('1','0','1','0','1','0','0','0','1','0','1','1','0','0'),
            ('1','0','1','0','1','0','0','0','1','0','1','1','1','0'),
            ('1','0','1','0','1','0','0','0','1','1','0','0','0','0'),
            ('1','0','1','0','1','0','0','0','1','1','0','0','1','0'),
            ('1','0','1','0','1','0','0','0','1','1','0','1','0','0'),
            ('1','0','1','0','1','0','0','0','1','1','0','1','1','0'),
            ('1','0','1','0','1','0','0','0','1','1','1','0','0','0'),
            ('1','0','1','0','1','0','0','0','1','1','1','0','1','0'),
            ('1','0','1','0','1','0','0','0','1','1','1','1','0','0'),
            ('1','0','1','0','1','0','0','0','1','1','1','1','1','0'),
            ('1','0','1','0','1','0','0','1','0','0','0','0','0','0'),
            ('1','0','1','0','1','0','0','1','0','0','0','0','1','0'),
            ('1','0','1','0','1','0','0','1','0','0','0','1','0','0'),
            ('1','0','1','0','1','0','0','1','0','0','0','1','1','0'),
            ('1','0','1','0','1','0','0','1','0','0','1','0','0','0'),
            ('1','0','1','0','1','0','0','1','0','0','1','0','1','0'),
            ('1','0','1','0','1','0','0','1','0','0','1','1','0','0'),
            ('1','0','1','0','1','0','0','1','0','0','1','1','1','0'),
            ('1','0','1','0','1','0','0','1','0','1','0','0','0','0'),
            ('1','0','1','0','1','0','0','1','0','1','0','0','1','0'),
            ('1','0','1','0','1','0','0','1','0','1','0','1','0','0'),
            ('1','0','1','0','1','0','0','1','0','1','0','1','1','0'),
            ('1','0','1','0','1','0','0','1','0','1','1','0','0','0'),
            ('1','0','1','0','1','0','0','1','0','1','1','0','1','0'),
            ('1','0','1','0','1','0','0','1','0','1','1','1','0','0'),
            ('1','0','1','0','1','0','0','1','0','1','1','1','1','0'),
            ('1','0','1','0','1','0','0','1','1','0','0','0','0','0'),
            ('1','0','1','0','1','0','0','1','1','0','0','0','1','0'),
            ('1','0','1','0','1','0','0','1','1','0','0','1','0','0'),
            ('1','0','1','0','1','0','0','1','1','0','0','1','1','0'),
            ('1','0','1','0','1','0','0','1','1','0','1','0','0','0'),
            ('1','0','1','0','1','0','0','1','1','0','1','0','1','0'),
            ('1','0','1','0','1','0','0','1','1','0','1','1','0','0'),
            ('1','0','1','0','1','0','0','1','1','0','1','1','1','0'),
            ('1','0','1','0','1','0','0','1','1','1','0','0','0','0'),
            ('1','0','1','0','1','0','0','1','1','1','0','0','1','0'),
            ('1','0','1','0','1','0','0','1','1','1','0','1','0','0'),
            ('1','0','1','0','1','0','0','1','1','1','0','1','1','0'),
            ('1','0','1','0','1','0','0','1','1','1','1','0','0','0'),
            ('1','0','1','0','1','0','0','1','1','1','1','0','1','0'),
            ('1','0','1','0','1','0','0','1','1','1','1','1','0','0'),
            ('1','0','1','0','1','0','0','1','1','1','1','1','1','0'),
            ('1','0','1','0','1','0','1','0','0','0','0','0','0','0'),
            ('1','0','1','0','1','0','1','0','0','0','0','0','1','0'),
            ('1','0','1','0','1','0','1','0','0','0','0','1','0','0'),
            ('1','0','1','0','1','0','1','0','0','0','0','1','1','0'),
            ('1','0','1','0','1','0','1','0','0','0','1','0','0','0'),
            ('1','0','1','0','1','0','1','0','0','0','1','0','1','0'),
            ('1','0','1','0','1','0','1','0','0','0','1','1','0','0'),
            ('1','0','1','0','1','0','1','0','0','0','1','1','1','0'),
            ('1','0','1','0','1','0','1','0','0','1','0','0','0','0'),
            ('1','0','1','0','1','0','1','0','0','1','0','0','1','0'),
            ('1','0','1','0','1','0','1','0','0','1','0','1','0','0'),
            ('1','0','1','0','1','0','1','0','0','1','0','1','1','0'),
            ('1','0','1','0','1','0','1','0','0','1','1','0','0','0'),
            ('1','0','1','0','1','0','1','0','0','1','1','0','1','0'),
            ('1','0','1','0','1','0','1','0','0','1','1','1','0','0'),
            ('1','0','1','0','1','0','1','0','0','1','1','1','1','0'),
            ('1','0','1','0','1','0','1','0','1','0','0','0','0','0'),
            ('1','0','1','0','1','0','1','0','1','0','0','0','1','0'),
            ('1','0','1','0','1','0','1','0','1','0','0','1','0','0'),
            ('1','0','1','0','1','0','1','0','1','0','0','1','1','0'),
            ('1','0','1','0','1','0','1','0','1','0','1','0','0','0'),
            ('1','0','1','0','1','0','1','0','1','0','1','0','1','0'),
            ('1','0','1','0','1','0','1','0','1','0','1','1','0','0'),
            ('1','0','1','0','1','0','1','0','1','0','1','1','1','0'),
            ('1','0','1','0','1','0','1','0','1','1','0','0','0','0'),
            ('1','0','1','0','1','0','1','0','1','1','0','0','1','0'),
            ('1','0','1','0','1','0','1','0','1','1','0','1','0','0'),
            ('1','0','1','0','1','0','1','0','1','1','0','1','1','0'),
            ('1','0','1','0','1','0','1','0','1','1','1','0','0','0'),
            ('1','0','1','0','1','0','1','0','1','1','1','0','1','0'),
            ('1','0','1','0','1','0','1','0','1','1','1','1','0','0'),
            ('1','0','1','0','1','0','1','0','1','1','1','1','1','0'),
            ('1','0','1','0','1','0','1','1','0','0','0','0','0','0'),
            ('1','0','1','0','1','0','1','1','0','0','0','0','1','0'),
            ('1','0','1','0','1','0','1','1','0','0','0','1','0','0'),
            ('1','0','1','0','1','0','1','1','0','0','0','1','1','0'),
            ('1','0','1','0','1','0','1','1','0','0','1','0','0','0'),
            ('1','0','1','0','1','0','1','1','0','0','1','0','1','0'),
            ('1','0','1','0','1','0','1','1','0','0','1','1','0','0'),
            ('1','0','1','0','1','0','1','1','0','0','1','1','1','0'),
            ('1','0','1','0','1','0','1','1','0','1','0','0','0','0'),
            ('1','0','1','0','1','0','1','1','0','1','0','0','1','0'),
            ('1','0','1','0','1','0','1','1','0','1','0','1','0','0'),
            ('1','0','1','0','1','0','1','1','0','1','0','1','1','0'),
            ('1','0','1','0','1','0','1','1','0','1','1','0','0','0'),
            ('1','0','1','0','1','0','1','1','0','1','1','0','1','0'),
            ('1','0','1','0','1','0','1','1','0','1','1','1','0','0'),
            ('1','0','1','0','1','0','1','1','0','1','1','1','1','0'),
            ('1','0','1','0','1','0','1','1','1','0','0','0','0','0'),
            ('1','0','1','0','1','0','1','1','1','0','0','0','1','0'),
            ('1','0','1','0','1','0','1','1','1','0','0','1','0','0'),
            ('1','0','1','0','1','0','1','1','1','0','0','1','1','0'),
            ('1','0','1','0','1','0','1','1','1','0','1','0','0','0'),
            ('1','0','1','0','1','0','1','1','1','0','1','0','1','0'),
            ('1','0','1','0','1','0','1','1','1','0','1','1','0','0'),
            ('1','0','1','0','1','0','1','1','1','0','1','1','1','0'),
            ('1','0','1','0','1','0','1','1','1','1','0','0','0','0'),
            ('1','0','1','0','1','0','1','1','1','1','0','0','1','0'),
            ('1','0','1','0','1','0','1','1','1','1','0','1','0','0'),
            ('1','0','1','0','1','0','1','1','1','1','0','1','1','0'),
            ('1','0','1','0','1','0','1','1','1','1','1','0','0','0'),
            ('1','0','1','0','1','0','1','1','1','1','1','0','1','0'),
            ('1','0','1','0','1','0','1','1','1','1','1','1','0','0'),
            ('1','0','1','0','1','0','1','1','1','1','1','1','1','0'),
            ('1','0','1','0','1','1','0','0','0','0','0','0','0','0'),
            ('1','0','1','0','1','1','0','0','0','0','0','0','1','0'),
            ('1','0','1','0','1','1','0','0','0','0','0','1','0','0'),
            ('1','0','1','0','1','1','0','0','0','0','0','1','1','0'),
            ('1','0','1','0','1','1','0','0','0','0','1','0','0','0'),
            ('1','0','1','0','1','1','0','0','0','0','1','0','1','0'),
            ('1','0','1','0','1','1','0','0','0','0','1','1','0','0'),
            ('1','0','1','0','1','1','0','0','0','0','1','1','1','0'),
            ('1','0','1','0','1','1','0','0','0','1','0','0','0','0'),
            ('1','0','1','0','1','1','0','0','0','1','0','0','1','0'),
            ('1','0','1','0','1','1','0','0','0','1','0','1','0','0'),
            ('1','0','1','0','1','1','0','0','0','1','0','1','1','0'),
            ('1','0','1','0','1','1','0','0','0','1','1','0','0','0'),
            ('1','0','1','0','1','1','0','0','0','1','1','0','1','0'),
            ('1','0','1','0','1','1','0','0','0','1','1','1','0','0'),
            ('1','0','1','0','1','1','0','0','0','1','1','1','1','0'),
            ('1','0','1','0','1','1','0','0','1','0','0','0','0','0'),
            ('1','0','1','0','1','1','0','0','1','0','0','0','1','0'),
            ('1','0','1','0','1','1','0','0','1','0','0','1','0','0'),
            ('1','0','1','0','1','1','0','0','1','0','0','1','1','0'),
            ('1','0','1','0','1','1','0','0','1','0','1','0','0','0'),
            ('1','0','1','0','1','1','0','0','1','0','1','0','1','0'),
            ('1','0','1','0','1','1','0','0','1','0','1','1','0','0'),
            ('1','0','1','0','1','1','0','0','1','0','1','1','1','0'),
            ('1','0','1','0','1','1','0','0','1','1','0','0','0','0'),
            ('1','0','1','0','1','1','0','0','1','1','0','0','1','0'),
            ('1','0','1','0','1','1','0','0','1','1','0','1','0','0'),
            ('1','0','1','0','1','1','0','0','1','1','0','1','1','0'),
            ('1','0','1','0','1','1','0','0','1','1','1','0','0','0'),
            ('1','0','1','0','1','1','0','0','1','1','1','0','1','0'),
            ('1','0','1','0','1','1','0','0','1','1','1','1','0','0'),
            ('1','0','1','0','1','1','0','0','1','1','1','1','1','0'),
            ('1','0','1','0','1','1','0','1','0','0','0','0','0','0'),
            ('1','0','1','0','1','1','0','1','0','0','0','0','1','0'),
            ('1','0','1','0','1','1','0','1','0','0','0','1','0','0'),
            ('1','0','1','0','1','1','0','1','0','0','0','1','1','0'),
            ('1','0','1','0','1','1','0','1','0','0','1','0','0','0'),
            ('1','0','1','0','1','1','0','1','0','0','1','0','1','0'),
            ('1','0','1','0','1','1','0','1','0','0','1','1','0','0'),
            ('1','0','1','0','1','1','0','1','0','0','1','1','1','0'),
            ('1','0','1','0','1','1','0','1','0','1','0','0','0','0'),
            ('1','0','1','0','1','1','0','1','0','1','0','0','1','0'),
            ('1','0','1','0','1','1','0','1','0','1','0','1','0','0'),
            ('1','0','1','0','1','1','0','1','0','1','0','1','1','0'),
            ('1','0','1','0','1','1','0','1','0','1','1','0','0','0'),
            ('1','0','1','0','1','1','0','1','0','1','1','0','1','0'),
            ('1','0','1','0','1','1','0','1','0','1','1','1','0','0'),
            ('1','0','1','0','1','1','0','1','0','1','1','1','1','0'),
            ('1','0','1','0','1','1','0','1','1','0','0','0','0','0'),
            ('1','0','1','0','1','1','0','1','1','0','0','0','1','0'),
            ('1','0','1','0','1','1','0','1','1','0','0','1','0','0'),
            ('1','0','1','0','1','1','0','1','1','0','0','1','1','0'),
            ('1','0','1','0','1','1','0','1','1','0','1','0','0','0'),
            ('1','0','1','0','1','1','0','1','1','0','1','0','1','0'),
            ('1','0','1','0','1','1','0','1','1','0','1','1','0','0'),
            ('1','0','1','0','1','1','0','1','1','0','1','1','1','0'),
            ('1','0','1','0','1','1','0','1','1','1','0','0','0','0'),
            ('1','0','1','0','1','1','0','1','1','1','0','0','1','0'),
            ('1','0','1','0','1','1','0','1','1','1','0','1','0','0'),
            ('1','0','1','0','1','1','0','1','1','1','0','1','1','0'),
            ('1','0','1','0','1','1','0','1','1','1','1','0','0','0'),
            ('1','0','1','0','1','1','0','1','1','1','1','0','1','0'),
            ('1','0','1','0','1','1','0','1','1','1','1','1','0','0'),
            ('1','0','1','0','1','1','0','1','1','1','1','1','1','0'),
            ('1','0','1','0','1','1','1','0','0','0','0','0','0','0'),
            ('1','0','1','0','1','1','1','0','0','0','0','0','1','0'),
            ('1','0','1','0','1','1','1','0','0','0','0','1','0','0'),
            ('1','0','1','0','1','1','1','0','0','0','0','1','1','0'),
            ('1','0','1','0','1','1','1','0','0','0','1','0','0','0'),
            ('1','0','1','0','1','1','1','0','0','0','1','0','1','0'),
            ('1','0','1','0','1','1','1','0','0','0','1','1','0','0'),
            ('1','0','1','0','1','1','1','0','0','0','1','1','1','0'),
            ('1','0','1','0','1','1','1','0','0','1','0','0','0','0'),
            ('1','0','1','0','1','1','1','0','0','1','0','0','1','0'),
            ('1','0','1','0','1','1','1','0','0','1','0','1','0','0'),
            ('1','0','1','0','1','1','1','0','0','1','0','1','1','0'),
            ('1','0','1','0','1','1','1','0','0','1','1','0','0','0'),
            ('1','0','1','0','1','1','1','0','0','1','1','0','1','0'),
            ('1','0','1','0','1','1','1','0','0','1','1','1','0','0'),
            ('1','0','1','0','1','1','1','0','0','1','1','1','1','0'),
            ('1','0','1','0','1','1','1','0','1','0','0','0','0','0'),
            ('1','0','1','0','1','1','1','0','1','0','0','0','1','0'),
            ('1','0','1','0','1','1','1','0','1','0','0','1','0','0'),
            ('1','0','1','0','1','1','1','0','1','0','0','1','1','0'),
            ('1','0','1','0','1','1','1','0','1','0','1','0','0','0'),
            ('1','0','1','0','1','1','1','0','1','0','1','0','1','0'),
            ('1','0','1','0','1','1','1','0','1','0','1','1','0','0'),
            ('1','0','1','0','1','1','1','0','1','0','1','1','1','0'),
            ('1','0','1','0','1','1','1','0','1','1','0','0','0','0'),
            ('1','0','1','0','1','1','1','0','1','1','0','0','1','0'),
            ('1','0','1','0','1','1','1','0','1','1','0','1','0','0'),
            ('1','0','1','0','1','1','1','0','1','1','0','1','1','0'),
            ('1','0','1','0','1','1','1','0','1','1','1','0','0','0'),
            ('1','0','1','0','1','1','1','0','1','1','1','0','1','0'),
            ('1','0','1','0','1','1','1','0','1','1','1','1','0','0'),
            ('1','0','1','0','1','1','1','0','1','1','1','1','1','0'),
            ('1','0','1','0','1','1','1','1','0','0','0','0','0','0'),
            ('1','0','1','0','1','1','1','1','0','0','0','0','1','0'),
            ('1','0','1','0','1','1','1','1','0','0','0','1','0','0'),
            ('1','0','1','0','1','1','1','1','0','0','0','1','1','0'),
            ('1','0','1','0','1','1','1','1','0','0','1','0','0','0'),
            ('1','0','1','0','1','1','1','1','0','0','1','0','1','0'),
            ('1','0','1','0','1','1','1','1','0','0','1','1','0','0'),
            ('1','0','1','0','1','1','1','1','0','0','1','1','1','0'),
            ('1','0','1','0','1','1','1','1','0','1','0','0','0','0'),
            ('1','0','1','0','1','1','1','1','0','1','0','0','1','0'),
            ('1','0','1','0','1','1','1','1','0','1','0','1','0','0'),
            ('1','0','1','0','1','1','1','1','0','1','0','1','1','0'),
            ('1','0','1','0','1','1','1','1','0','1','1','0','0','0'),
            ('1','0','1','0','1','1','1','1','0','1','1','0','1','0'),
            ('1','0','1','0','1','1','1','1','0','1','1','1','0','0'),
            ('1','0','1','0','1','1','1','1','0','1','1','1','1','0'),
            ('1','0','1','0','1','1','1','1','1','0','0','0','0','0'),
            ('1','0','1','0','1','1','1','1','1','0','0','0','1','0'),
            ('1','0','1','0','1','1','1','1','1','0','0','1','0','0'),
            ('1','0','1','0','1','1','1','1','1','0','0','1','1','0'),
            ('1','0','1','0','1','1','1','1','1','0','1','0','0','0'),
            ('1','0','1','0','1','1','1','1','1','0','1','0','1','0'),
            ('1','0','1','0','1','1','1','1','1','0','1','1','0','0'),
            ('1','0','1','0','1','1','1','1','1','0','1','1','1','0'),
            ('1','0','1','0','1','1','1','1','1','1','0','0','0','0'),
            ('1','0','1','0','1','1','1','1','1','1','0','0','1','0'),
            ('1','0','1','0','1','1','1','1','1','1','0','1','0','0'),
            ('1','0','1','0','1','1','1','1','1','1','0','1','1','0'),
            ('1','0','1','0','1','1','1','1','1','1','1','0','0','0'),
            ('1','0','1','0','1','1','1','1','1','1','1','0','1','0'),
            ('1','0','1','0','1','1','1','1','1','1','1','1','0','0'),
            ('1','0','1','0','1','1','1','1','1','1','1','1','1','0'),
            ('1','0','1','1','0','0','0','0','0','0','0','0','0','0'),
            ('1','0','1','1','0','0','0','0','0','0','0','0','1','0'),
            ('1','0','1','1','0','0','0','0','0','0','0','1','0','0'),
            ('1','0','1','1','0','0','0','0','0','0','0','1','1','0'),
            ('1','0','1','1','0','0','0','0','0','0','1','0','0','0'),
            ('1','0','1','1','0','0','0','0','0','0','1','0','1','0'),
            ('1','0','1','1','0','0','0','0','0','0','1','1','0','0'),
            ('1','0','1','1','0','0','0','0','0','0','1','1','1','0'),
            ('1','0','1','1','0','0','0','0','0','1','0','0','0','0'),
            ('1','0','1','1','0','0','0','0','0','1','0','0','1','0'),
            ('1','0','1','1','0','0','0','0','0','1','0','1','0','0'),
            ('1','0','1','1','0','0','0','0','0','1','0','1','1','0'),
            ('1','0','1','1','0','0','0','0','0','1','1','0','0','0'),
            ('1','0','1','1','0','0','0','0','0','1','1','0','1','0'),
            ('1','0','1','1','0','0','0','0','0','1','1','1','0','0'),
            ('1','0','1','1','0','0','0','0','0','1','1','1','1','0'),
            ('1','0','1','1','0','0','0','0','1','0','0','0','0','0'),
            ('1','0','1','1','0','0','0','0','1','0','0','0','1','0'),
            ('1','0','1','1','0','0','0','0','1','0','0','1','0','0'),
            ('1','0','1','1','0','0','0','0','1','0','0','1','1','0'),
            ('1','0','1','1','0','0','0','0','1','0','1','0','0','0'),
            ('1','0','1','1','0','0','0','0','1','0','1','0','1','0'),
            ('1','0','1','1','0','0','0','0','1','0','1','1','0','0'),
            ('1','0','1','1','0','0','0','0','1','0','1','1','1','0'),
            ('1','0','1','1','0','0','0','0','1','1','0','0','0','0'),
            ('1','0','1','1','0','0','0','0','1','1','0','0','1','0'),
            ('1','0','1','1','0','0','0','0','1','1','0','1','0','0'),
            ('1','0','1','1','0','0','0','0','1','1','0','1','1','0'),
            ('1','0','1','1','0','0','0','0','1','1','1','0','0','0'),
            ('1','0','1','1','0','0','0','0','1','1','1','0','1','0'),
            ('1','0','1','1','0','0','0','0','1','1','1','1','0','0'),
            ('1','0','1','1','0','0','0','0','1','1','1','1','1','0'),
            ('1','0','1','1','0','0','0','1','0','0','0','0','0','0'),
            ('1','0','1','1','0','0','0','1','0','0','0','0','1','0'),
            ('1','0','1','1','0','0','0','1','0','0','0','1','0','0'),
            ('1','0','1','1','0','0','0','1','0','0','0','1','1','0'),
            ('1','0','1','1','0','0','0','1','0','0','1','0','0','0'),
            ('1','0','1','1','0','0','0','1','0','0','1','0','1','0'),
            ('1','0','1','1','0','0','0','1','0','0','1','1','0','0'),
            ('1','0','1','1','0','0','0','1','0','0','1','1','1','0'),
            ('1','0','1','1','0','0','0','1','0','1','0','0','0','0'),
            ('1','0','1','1','0','0','0','1','0','1','0','0','1','0'),
            ('1','0','1','1','0','0','0','1','0','1','0','1','0','0'),
            ('1','0','1','1','0','0','0','1','0','1','0','1','1','0'),
            ('1','0','1','1','0','0','0','1','0','1','1','0','0','0'),
            ('1','0','1','1','0','0','0','1','0','1','1','0','1','0'),
            ('1','0','1','1','0','0','0','1','0','1','1','1','0','0'),
            ('1','0','1','1','0','0','0','1','0','1','1','1','1','0'),
            ('1','0','1','1','0','0','0','1','1','0','0','0','0','0'),
            ('1','0','1','1','0','0','0','1','1','0','0','0','1','0'),
            ('1','0','1','1','0','0','0','1','1','0','0','1','0','0'),
            ('1','0','1','1','0','0','0','1','1','0','0','1','1','0'),
            ('1','0','1','1','0','0','0','1','1','0','1','0','0','0'),
            ('1','0','1','1','0','0','0','1','1','0','1','0','1','0'),
            ('1','0','1','1','0','0','0','1','1','0','1','1','0','0'),
            ('1','0','1','1','0','0','0','1','1','0','1','1','1','0'),
            ('1','0','1','1','0','0','0','1','1','1','0','0','0','0'),
            ('1','0','1','1','0','0','0','1','1','1','0','0','1','0'),
            ('1','0','1','1','0','0','0','1','1','1','0','1','0','0'),
            ('1','0','1','1','0','0','0','1','1','1','0','1','1','0'),
            ('1','0','1','1','0','0','0','1','1','1','1','0','0','0'),
            ('1','0','1','1','0','0','0','1','1','1','1','0','1','0'),
            ('1','0','1','1','0','0','0','1','1','1','1','1','0','0'),
            ('1','0','1','1','0','0','0','1','1','1','1','1','1','0'),
            ('1','0','1','1','0','0','1','0','0','0','0','0','0','0'),
            ('1','0','1','1','0','0','1','0','0','0','0','0','1','0'),
            ('1','0','1','1','0','0','1','0','0','0','0','1','0','0'),
            ('1','0','1','1','0','0','1','0','0','0','0','1','1','0'),
            ('1','0','1','1','0','0','1','0','0','0','1','0','0','0'),
            ('1','0','1','1','0','0','1','0','0','0','1','0','1','0'),
            ('1','0','1','1','0','0','1','0','0','0','1','1','0','0'),
            ('1','0','1','1','0','0','1','0','0','0','1','1','1','0'),
            ('1','0','1','1','0','0','1','0','0','1','0','0','0','0'),
            ('1','0','1','1','0','0','1','0','0','1','0','0','1','0'),
            ('1','0','1','1','0','0','1','0','0','1','0','1','0','0'),
            ('1','0','1','1','0','0','1','0','0','1','0','1','1','0'),
            ('1','0','1','1','0','0','1','0','0','1','1','0','0','0'),
            ('1','0','1','1','0','0','1','0','0','1','1','0','1','0'),
            ('1','0','1','1','0','0','1','0','0','1','1','1','0','0'),
            ('1','0','1','1','0','0','1','0','0','1','1','1','1','0'),
            ('1','0','1','1','0','0','1','0','1','0','0','0','0','0'),
            ('1','0','1','1','0','0','1','0','1','0','0','0','1','0'),
            ('1','0','1','1','0','0','1','0','1','0','0','1','0','0'),
            ('1','0','1','1','0','0','1','0','1','0','0','1','1','0'),
            ('1','0','1','1','0','0','1','0','1','0','1','0','0','0'),
            ('1','0','1','1','0','0','1','0','1','0','1','0','1','0'),
            ('1','0','1','1','0','0','1','0','1','0','1','1','0','0'),
            ('1','0','1','1','0','0','1','0','1','0','1','1','1','0'),
            ('1','0','1','1','0','0','1','0','1','1','0','0','0','0'),
            ('1','0','1','1','0','0','1','0','1','1','0','0','1','0'),
            ('1','0','1','1','0','0','1','0','1','1','0','1','0','0'),
            ('1','0','1','1','0','0','1','0','1','1','0','1','1','0'),
            ('1','0','1','1','0','0','1','0','1','1','1','0','0','0'),
            ('1','0','1','1','0','0','1','0','1','1','1','0','1','0'),
            ('1','0','1','1','0','0','1','0','1','1','1','1','0','0'),
            ('1','0','1','1','0','0','1','0','1','1','1','1','1','0'),
            ('1','0','1','1','0','0','1','1','0','0','0','0','0','0'),
            ('1','0','1','1','0','0','1','1','0','0','0','0','1','0'),
            ('1','0','1','1','0','0','1','1','0','0','0','1','0','0'),
            ('1','0','1','1','0','0','1','1','0','0','0','1','1','0'),
            ('1','0','1','1','0','0','1','1','0','0','1','0','0','0'),
            ('1','0','1','1','0','0','1','1','0','0','1','0','1','0'),
            ('1','0','1','1','0','0','1','1','0','0','1','1','0','0'),
            ('1','0','1','1','0','0','1','1','0','0','1','1','1','0'),
            ('1','0','1','1','0','0','1','1','0','1','0','0','0','0'),
            ('1','0','1','1','0','0','1','1','0','1','0','0','1','0'),
            ('1','0','1','1','0','0','1','1','0','1','0','1','0','0'),
            ('1','0','1','1','0','0','1','1','0','1','0','1','1','0'),
            ('1','0','1','1','0','0','1','1','0','1','1','0','0','0'),
            ('1','0','1','1','0','0','1','1','0','1','1','0','1','0'),
            ('1','0','1','1','0','0','1','1','0','1','1','1','0','0'),
            ('1','0','1','1','0','0','1','1','0','1','1','1','1','0'),
            ('1','0','1','1','0','0','1','1','1','0','0','0','0','0'),
            ('1','0','1','1','0','0','1','1','1','0','0','0','1','0'),
            ('1','0','1','1','0','0','1','1','1','0','0','1','0','0'),
            ('1','0','1','1','0','0','1','1','1','0','0','1','1','0'),
            ('1','0','1','1','0','0','1','1','1','0','1','0','0','0'),
            ('1','0','1','1','0','0','1','1','1','0','1','0','1','0'),
            ('1','0','1','1','0','0','1','1','1','0','1','1','0','0'),
            ('1','0','1','1','0','0','1','1','1','0','1','1','1','0'),
            ('1','0','1','1','0','0','1','1','1','1','0','0','0','0'),
            ('1','0','1','1','0','0','1','1','1','1','0','0','1','0'),
            ('1','0','1','1','0','0','1','1','1','1','0','1','0','0'),
            ('1','0','1','1','0','0','1','1','1','1','0','1','1','0'),
            ('1','0','1','1','0','0','1','1','1','1','1','0','0','0'),
            ('1','0','1','1','0','0','1','1','1','1','1','0','1','0'),
            ('1','0','1','1','0','0','1','1','1','1','1','1','0','0'),
            ('1','0','1','1','0','0','1','1','1','1','1','1','1','0'),
            ('1','0','1','1','0','1','0','0','0','0','0','0','0','0'),
            ('1','0','1','1','0','1','0','0','0','0','0','0','1','0'),
            ('1','0','1','1','0','1','0','0','0','0','0','1','0','0'),
            ('1','0','1','1','0','1','0','0','0','0','0','1','1','0'),
            ('1','0','1','1','0','1','0','0','0','0','1','0','0','0'),
            ('1','0','1','1','0','1','0','0','0','0','1','0','1','0'),
            ('1','0','1','1','0','1','0','0','0','0','1','1','0','0'),
            ('1','0','1','1','0','1','0','0','0','0','1','1','1','0'),
            ('1','0','1','1','0','1','0','0','0','1','0','0','0','0'),
            ('1','0','1','1','0','1','0','0','0','1','0','0','1','0'),
            ('1','0','1','1','0','1','0','0','0','1','0','1','0','0'),
            ('1','0','1','1','0','1','0','0','0','1','0','1','1','0'),
            ('1','0','1','1','0','1','0','0','0','1','1','0','0','0'),
            ('1','0','1','1','0','1','0','0','0','1','1','0','1','0'),
            ('1','0','1','1','0','1','0','0','0','1','1','1','0','0'),
            ('1','0','1','1','0','1','0','0','0','1','1','1','1','0'),
            ('1','0','1','1','0','1','0','0','1','0','0','0','0','0'),
            ('1','0','1','1','0','1','0','0','1','0','0','0','1','0'),
            ('1','0','1','1','0','1','0','0','1','0','0','1','0','0'),
            ('1','0','1','1','0','1','0','0','1','0','0','1','1','0'),
            ('1','0','1','1','0','1','0','0','1','0','1','0','0','0'),
            ('1','0','1','1','0','1','0','0','1','0','1','0','1','0'),
            ('1','0','1','1','0','1','0','0','1','0','1','1','0','0'),
            ('1','0','1','1','0','1','0','0','1','0','1','1','1','0'),
            ('1','0','1','1','0','1','0','0','1','1','0','0','0','0'),
            ('1','0','1','1','0','1','0','0','1','1','0','0','1','0'),
            ('1','0','1','1','0','1','0','0','1','1','0','1','0','0'),
            ('1','0','1','1','0','1','0','0','1','1','0','1','1','0'),
            ('1','0','1','1','0','1','0','0','1','1','1','0','0','0'),
            ('1','0','1','1','0','1','0','0','1','1','1','0','1','0'),
            ('1','0','1','1','0','1','0','0','1','1','1','1','0','0'),
            ('1','0','1','1','0','1','0','0','1','1','1','1','1','0'),
            ('1','0','1','1','0','1','0','1','0','0','0','0','0','0'),
            ('1','0','1','1','0','1','0','1','0','0','0','0','1','0'),
            ('1','0','1','1','0','1','0','1','0','0','0','1','0','0'),
            ('1','0','1','1','0','1','0','1','0','0','0','1','1','0'),
            ('1','0','1','1','0','1','0','1','0','0','1','0','0','0'),
            ('1','0','1','1','0','1','0','1','0','0','1','0','1','0'),
            ('1','0','1','1','0','1','0','1','0','0','1','1','0','0'),
            ('1','0','1','1','0','1','0','1','0','0','1','1','1','0'),
            ('1','0','1','1','0','1','0','1','0','1','0','0','0','0'),
            ('1','0','1','1','0','1','0','1','0','1','0','0','1','0'),
            ('1','0','1','1','0','1','0','1','0','1','0','1','0','0'),
            ('1','0','1','1','0','1','0','1','0','1','0','1','1','0'),
            ('1','0','1','1','0','1','0','1','0','1','1','0','0','0'),
            ('1','0','1','1','0','1','0','1','0','1','1','0','1','0'),
            ('1','0','1','1','0','1','0','1','0','1','1','1','0','0'),
            ('1','0','1','1','0','1','0','1','0','1','1','1','1','0'),
            ('1','0','1','1','0','1','0','1','1','0','0','0','0','0'),
            ('1','0','1','1','0','1','0','1','1','0','0','0','1','0'),
            ('1','0','1','1','0','1','0','1','1','0','0','1','0','0'),
            ('1','0','1','1','0','1','0','1','1','0','0','1','1','0'),
            ('1','0','1','1','0','1','0','1','1','0','1','0','0','0'),
            ('1','0','1','1','0','1','0','1','1','0','1','0','1','0'),
            ('1','0','1','1','0','1','0','1','1','0','1','1','0','0'),
            ('1','0','1','1','0','1','0','1','1','0','1','1','1','0'),
            ('1','0','1','1','0','1','0','1','1','1','0','0','0','0'),
            ('1','0','1','1','0','1','0','1','1','1','0','0','1','0'),
            ('1','0','1','1','0','1','0','1','1','1','0','1','0','0'),
            ('1','0','1','1','0','1','0','1','1','1','0','1','1','0'),
            ('1','0','1','1','0','1','0','1','1','1','1','0','0','0'),
            ('1','0','1','1','0','1','0','1','1','1','1','0','1','0'),
            ('1','0','1','1','0','1','0','1','1','1','1','1','0','0'),
            ('1','0','1','1','0','1','0','1','1','1','1','1','1','0'),
            ('1','0','1','1','0','1','1','0','0','0','0','0','0','0'),
            ('1','0','1','1','0','1','1','0','0','0','0','0','1','0'),
            ('1','0','1','1','0','1','1','0','0','0','0','1','0','0'),
            ('1','0','1','1','0','1','1','0','0','0','0','1','1','0'),
            ('1','0','1','1','0','1','1','0','0','0','1','0','0','0'),
            ('1','0','1','1','0','1','1','0','0','0','1','0','1','0'),
            ('1','0','1','1','0','1','1','0','0','0','1','1','0','0'),
            ('1','0','1','1','0','1','1','0','0','0','1','1','1','0'),
            ('1','0','1','1','0','1','1','0','0','1','0','0','0','0'),
            ('1','0','1','1','0','1','1','0','0','1','0','0','1','0'),
            ('1','0','1','1','0','1','1','0','0','1','0','1','0','0'),
            ('1','0','1','1','0','1','1','0','0','1','0','1','1','0'),
            ('1','0','1','1','0','1','1','0','0','1','1','0','0','0'),
            ('1','0','1','1','0','1','1','0','0','1','1','0','1','0'),
            ('1','0','1','1','0','1','1','0','0','1','1','1','0','0'),
            ('1','0','1','1','0','1','1','0','0','1','1','1','1','0'),
            ('1','0','1','1','0','1','1','0','1','0','0','0','0','0'),
            ('1','0','1','1','0','1','1','0','1','0','0','0','1','0'),
            ('1','0','1','1','0','1','1','0','1','0','0','1','0','0'),
            ('1','0','1','1','0','1','1','0','1','0','0','1','1','0'),
            ('1','0','1','1','0','1','1','0','1','0','1','0','0','0'),
            ('1','0','1','1','0','1','1','0','1','0','1','0','1','0'),
            ('1','0','1','1','0','1','1','0','1','0','1','1','0','0'),
            ('1','0','1','1','0','1','1','0','1','0','1','1','1','0'),
            ('1','0','1','1','0','1','1','0','1','1','0','0','0','0'),
            ('1','0','1','1','0','1','1','0','1','1','0','0','1','0'),
            ('1','0','1','1','0','1','1','0','1','1','0','1','0','0'),
            ('1','0','1','1','0','1','1','0','1','1','0','1','1','0'),
            ('1','0','1','1','0','1','1','0','1','1','1','0','0','0'),
            ('1','0','1','1','0','1','1','0','1','1','1','0','1','0'),
            ('1','0','1','1','0','1','1','0','1','1','1','1','0','0'),
            ('1','0','1','1','0','1','1','0','1','1','1','1','1','0'),
            ('1','0','1','1','0','1','1','1','0','0','0','0','0','0'),
            ('1','0','1','1','0','1','1','1','0','0','0','0','1','0'),
            ('1','0','1','1','0','1','1','1','0','0','0','1','0','0'),
            ('1','0','1','1','0','1','1','1','0','0','0','1','1','0'),
            ('1','0','1','1','0','1','1','1','0','0','1','0','0','0'),
            ('1','0','1','1','0','1','1','1','0','0','1','0','1','0'),
            ('1','0','1','1','0','1','1','1','0','0','1','1','0','0'),
            ('1','0','1','1','0','1','1','1','0','0','1','1','1','0'),
            ('1','0','1','1','0','1','1','1','0','1','0','0','0','0'),
            ('1','0','1','1','0','1','1','1','0','1','0','0','1','0'),
            ('1','0','1','1','0','1','1','1','0','1','0','1','0','0'),
            ('1','0','1','1','0','1','1','1','0','1','0','1','1','0'),
            ('1','0','1','1','0','1','1','1','0','1','1','0','0','0'),
            ('1','0','1','1','0','1','1','1','0','1','1','0','1','0'),
            ('1','0','1','1','0','1','1','1','0','1','1','1','0','0'),
            ('1','0','1','1','0','1','1','1','0','1','1','1','1','0'),
            ('1','0','1','1','0','1','1','1','1','0','0','0','0','0'),
            ('1','0','1','1','0','1','1','1','1','0','0','0','1','0'),
            ('1','0','1','1','0','1','1','1','1','0','0','1','0','0'),
            ('1','0','1','1','0','1','1','1','1','0','0','1','1','0'),
            ('1','0','1','1','0','1','1','1','1','0','1','0','0','0'),
            ('1','0','1','1','0','1','1','1','1','0','1','0','1','0'),
            ('1','0','1','1','0','1','1','1','1','0','1','1','0','0'),
            ('1','0','1','1','0','1','1','1','1','0','1','1','1','0'),
            ('1','0','1','1','0','1','1','1','1','1','0','0','0','0'),
            ('1','0','1','1','0','1','1','1','1','1','0','0','1','0'),
            ('1','0','1','1','0','1','1','1','1','1','0','1','0','0'),
            ('1','0','1','1','0','1','1','1','1','1','0','1','1','0'),
            ('1','0','1','1','0','1','1','1','1','1','1','0','0','0'),
            ('1','0','1','1','0','1','1','1','1','1','1','0','1','0'),
            ('1','0','1','1','0','1','1','1','1','1','1','1','0','0'),
            ('1','0','1','1','0','1','1','1','1','1','1','1','1','0'),
            ('1','0','1','1','1','0','0','0','0','0','0','0','0','0'),
            ('1','0','1','1','1','0','0','0','0','0','0','0','1','0'),
            ('1','0','1','1','1','0','0','0','0','0','0','1','0','0'),
            ('1','0','1','1','1','0','0','0','0','0','0','1','1','0'),
            ('1','0','1','1','1','0','0','0','0','0','1','0','0','0'),
            ('1','0','1','1','1','0','0','0','0','0','1','0','1','0'),
            ('1','0','1','1','1','0','0','0','0','0','1','1','0','0'),
            ('1','0','1','1','1','0','0','0','0','0','1','1','1','0'),
            ('1','0','1','1','1','0','0','0','0','1','0','0','0','0'),
            ('1','0','1','1','1','0','0','0','0','1','0','0','1','0'),
            ('1','0','1','1','1','0','0','0','0','1','0','1','0','0'),
            ('1','0','1','1','1','0','0','0','0','1','0','1','1','0'),
            ('1','0','1','1','1','0','0','0','0','1','1','0','0','0'),
            ('1','0','1','1','1','0','0','0','0','1','1','0','1','0'),
            ('1','0','1','1','1','0','0','0','0','1','1','1','0','0'),
            ('1','0','1','1','1','0','0','0','0','1','1','1','1','0'),
            ('1','0','1','1','1','0','0','0','1','0','0','0','0','0'),
            ('1','0','1','1','1','0','0','0','1','0','0','0','1','0'),
            ('1','0','1','1','1','0','0','0','1','0','0','1','0','0'),
            ('1','0','1','1','1','0','0','0','1','0','0','1','1','0'),
            ('1','0','1','1','1','0','0','0','1','0','1','0','0','0'),
            ('1','0','1','1','1','0','0','0','1','0','1','0','1','0'),
            ('1','0','1','1','1','0','0','0','1','0','1','1','0','0'),
            ('1','0','1','1','1','0','0','0','1','0','1','1','1','0'),
            ('1','0','1','1','1','0','0','0','1','1','0','0','0','0'),
            ('1','0','1','1','1','0','0','0','1','1','0','0','1','0'),
            ('1','0','1','1','1','0','0','0','1','1','0','1','0','0'),
            ('1','0','1','1','1','0','0','0','1','1','0','1','1','0'),
            ('1','0','1','1','1','0','0','0','1','1','1','0','0','0'),
            ('1','0','1','1','1','0','0','0','1','1','1','0','1','0'),
            ('1','0','1','1','1','0','0','0','1','1','1','1','0','0'),
            ('1','0','1','1','1','0','0','0','1','1','1','1','1','0'),
            ('1','0','1','1','1','0','0','1','0','0','0','0','0','0'),
            ('1','0','1','1','1','0','0','1','0','0','0','0','1','0'),
            ('1','0','1','1','1','0','0','1','0','0','0','1','0','0'),
            ('1','0','1','1','1','0','0','1','0','0','0','1','1','0'),
            ('1','0','1','1','1','0','0','1','0','0','1','0','0','0'),
            ('1','0','1','1','1','0','0','1','0','0','1','0','1','0'),
            ('1','0','1','1','1','0','0','1','0','0','1','1','0','0'),
            ('1','0','1','1','1','0','0','1','0','0','1','1','1','0'),
            ('1','0','1','1','1','0','0','1','0','1','0','0','0','0'),
            ('1','0','1','1','1','0','0','1','0','1','0','0','1','0'),
            ('1','0','1','1','1','0','0','1','0','1','0','1','0','0'),
            ('1','0','1','1','1','0','0','1','0','1','0','1','1','0'),
            ('1','0','1','1','1','0','0','1','0','1','1','0','0','0'),
            ('1','0','1','1','1','0','0','1','0','1','1','0','1','0'),
            ('1','0','1','1','1','0','0','1','0','1','1','1','0','0'),
            ('1','0','1','1','1','0','0','1','0','1','1','1','1','0'),
            ('1','0','1','1','1','0','0','1','1','0','0','0','0','0'),
            ('1','0','1','1','1','0','0','1','1','0','0','0','1','0'),
            ('1','0','1','1','1','0','0','1','1','0','0','1','0','0'),
            ('1','0','1','1','1','0','0','1','1','0','0','1','1','0'),
            ('1','0','1','1','1','0','0','1','1','0','1','0','0','0'),
            ('1','0','1','1','1','0','0','1','1','0','1','0','1','0'),
            ('1','0','1','1','1','0','0','1','1','0','1','1','0','0'),
            ('1','0','1','1','1','0','0','1','1','0','1','1','1','0'),
            ('1','0','1','1','1','0','0','1','1','1','0','0','0','0'),
            ('1','0','1','1','1','0','0','1','1','1','0','0','1','0'),
            ('1','0','1','1','1','0','0','1','1','1','0','1','0','0'),
            ('1','0','1','1','1','0','0','1','1','1','0','1','1','0'),
            ('1','0','1','1','1','0','0','1','1','1','1','0','0','0'),
            ('1','0','1','1','1','0','0','1','1','1','1','0','1','0'),
            ('1','0','1','1','1','0','0','1','1','1','1','1','0','0'),
            ('1','0','1','1','1','0','0','1','1','1','1','1','1','0'),
            ('1','0','1','1','1','0','1','0','0','0','0','0','0','0'),
            ('1','0','1','1','1','0','1','0','0','0','0','0','1','0'),
            ('1','0','1','1','1','0','1','0','0','0','0','1','0','0'),
            ('1','0','1','1','1','0','1','0','0','0','0','1','1','0'),
            ('1','0','1','1','1','0','1','0','0','0','1','0','0','0'),
            ('1','0','1','1','1','0','1','0','0','0','1','0','1','0'),
            ('1','0','1','1','1','0','1','0','0','0','1','1','0','0'),
            ('1','0','1','1','1','0','1','0','0','0','1','1','1','0'),
            ('1','0','1','1','1','0','1','0','0','1','0','0','0','0'),
            ('1','0','1','1','1','0','1','0','0','1','0','0','1','0'),
            ('1','0','1','1','1','0','1','0','0','1','0','1','0','0'),
            ('1','0','1','1','1','0','1','0','0','1','0','1','1','0'),
            ('1','0','1','1','1','0','1','0','0','1','1','0','0','0'),
            ('1','0','1','1','1','0','1','0','0','1','1','0','1','0'),
            ('1','0','1','1','1','0','1','0','0','1','1','1','0','0'),
            ('1','0','1','1','1','0','1','0','0','1','1','1','1','0'),
            ('1','0','1','1','1','0','1','0','1','0','0','0','0','0'),
            ('1','0','1','1','1','0','1','0','1','0','0','0','1','0'),
            ('1','0','1','1','1','0','1','0','1','0','0','1','0','0'),
            ('1','0','1','1','1','0','1','0','1','0','0','1','1','0'),
            ('1','0','1','1','1','0','1','0','1','0','1','0','0','0'),
            ('1','0','1','1','1','0','1','0','1','0','1','0','1','0'),
            ('1','0','1','1','1','0','1','0','1','0','1','1','0','0'),
            ('1','0','1','1','1','0','1','0','1','0','1','1','1','0'),
            ('1','0','1','1','1','0','1','0','1','1','0','0','0','0'),
            ('1','0','1','1','1','0','1','0','1','1','0','0','1','0'),
            ('1','0','1','1','1','0','1','0','1','1','0','1','0','0'),
            ('1','0','1','1','1','0','1','0','1','1','0','1','1','0'),
            ('1','0','1','1','1','0','1','0','1','1','1','0','0','0'),
            ('1','0','1','1','1','0','1','0','1','1','1','0','1','0'),
            ('1','0','1','1','1','0','1','0','1','1','1','1','0','0'),
            ('1','0','1','1','1','0','1','0','1','1','1','1','1','0'),
            ('1','0','1','1','1','0','1','1','0','0','0','0','0','0'),
            ('1','0','1','1','1','0','1','1','0','0','0','0','1','0'),
            ('1','0','1','1','1','0','1','1','0','0','0','1','0','0'),
            ('1','0','1','1','1','0','1','1','0','0','0','1','1','0'),
            ('1','0','1','1','1','0','1','1','0','0','1','0','0','0'),
            ('1','0','1','1','1','0','1','1','0','0','1','0','1','0'),
            ('1','0','1','1','1','0','1','1','0','0','1','1','0','0'),
            ('1','0','1','1','1','0','1','1','0','0','1','1','1','0'),
            ('1','0','1','1','1','0','1','1','0','1','0','0','0','0'),
            ('1','0','1','1','1','0','1','1','0','1','0','0','1','0'),
            ('1','0','1','1','1','0','1','1','0','1','0','1','0','0'),
            ('1','0','1','1','1','0','1','1','0','1','0','1','1','0'),
            ('1','0','1','1','1','0','1','1','0','1','1','0','0','0'),
            ('1','0','1','1','1','0','1','1','0','1','1','0','1','0'),
            ('1','0','1','1','1','0','1','1','0','1','1','1','0','0'),
            ('1','0','1','1','1','0','1','1','0','1','1','1','1','0'),
            ('1','0','1','1','1','0','1','1','1','0','0','0','0','0'),
            ('1','0','1','1','1','0','1','1','1','0','0','0','1','0'),
            ('1','0','1','1','1','0','1','1','1','0','0','1','0','0'),
            ('1','0','1','1','1','0','1','1','1','0','0','1','1','0'),
            ('1','0','1','1','1','0','1','1','1','0','1','0','0','0'),
            ('1','0','1','1','1','0','1','1','1','0','1','0','1','0'),
            ('1','0','1','1','1','0','1','1','1','0','1','1','0','0'),
            ('1','0','1','1','1','0','1','1','1','0','1','1','1','0'),
            ('1','0','1','1','1','0','1','1','1','1','0','0','0','0'),
            ('1','0','1','1','1','0','1','1','1','1','0','0','1','0'),
            ('1','0','1','1','1','0','1','1','1','1','0','1','0','0'),
            ('1','0','1','1','1','0','1','1','1','1','0','1','1','0'),
            ('1','0','1','1','1','0','1','1','1','1','1','0','0','0'),
            ('1','0','1','1','1','0','1','1','1','1','1','0','1','0'),
            ('1','0','1','1','1','0','1','1','1','1','1','1','0','0'),
            ('1','0','1','1','1','0','1','1','1','1','1','1','1','0'),
            ('1','0','1','1','1','1','0','0','0','0','0','0','0','0'),
            ('1','0','1','1','1','1','0','0','0','0','0','0','1','0'),
            ('1','0','1','1','1','1','0','0','0','0','0','1','0','0'),
            ('1','0','1','1','1','1','0','0','0','0','0','1','1','0'),
            ('1','0','1','1','1','1','0','0','0','0','1','0','0','0'),
            ('1','0','1','1','1','1','0','0','0','0','1','0','1','0'),
            ('1','0','1','1','1','1','0','0','0','0','1','1','0','0'),
            ('1','0','1','1','1','1','0','0','0','0','1','1','1','0'),
            ('1','0','1','1','1','1','0','0','0','1','0','0','0','0'),
            ('1','0','1','1','1','1','0','0','0','1','0','0','1','0'),
            ('1','0','1','1','1','1','0','0','0','1','0','1','0','0'),
            ('1','0','1','1','1','1','0','0','0','1','0','1','1','0'),
            ('1','0','1','1','1','1','0','0','0','1','1','0','0','0'),
            ('1','0','1','1','1','1','0','0','0','1','1','0','1','0'),
            ('1','0','1','1','1','1','0','0','0','1','1','1','0','0'),
            ('1','0','1','1','1','1','0','0','0','1','1','1','1','0'),
            ('1','0','1','1','1','1','0','0','1','0','0','0','0','0'),
            ('1','0','1','1','1','1','0','0','1','0','0','0','1','0'),
            ('1','0','1','1','1','1','0','0','1','0','0','1','0','0'),
            ('1','0','1','1','1','1','0','0','1','0','0','1','1','0'),
            ('1','0','1','1','1','1','0','0','1','0','1','0','0','0'),
            ('1','0','1','1','1','1','0','0','1','0','1','0','1','0'),
            ('1','0','1','1','1','1','0','0','1','0','1','1','0','0'),
            ('1','0','1','1','1','1','0','0','1','0','1','1','1','0'),
            ('1','0','1','1','1','1','0','0','1','1','0','0','0','0'),
            ('1','0','1','1','1','1','0','0','1','1','0','0','1','0'),
            ('1','0','1','1','1','1','0','0','1','1','0','1','0','0'),
            ('1','0','1','1','1','1','0','0','1','1','0','1','1','0'),
            ('1','0','1','1','1','1','0','0','1','1','1','0','0','0'),
            ('1','0','1','1','1','1','0','0','1','1','1','0','1','0'),
            ('1','0','1','1','1','1','0','0','1','1','1','1','0','0'),
            ('1','0','1','1','1','1','0','0','1','1','1','1','1','0'),
            ('1','0','1','1','1','1','0','1','0','0','0','0','0','0'),
            ('1','0','1','1','1','1','0','1','0','0','0','0','1','0'),
            ('1','0','1','1','1','1','0','1','0','0','0','1','0','0'),
            ('1','0','1','1','1','1','0','1','0','0','0','1','1','0'),
            ('1','0','1','1','1','1','0','1','0','0','1','0','0','0'),
            ('1','0','1','1','1','1','0','1','0','0','1','0','1','0'),
            ('1','0','1','1','1','1','0','1','0','0','1','1','0','0'),
            ('1','0','1','1','1','1','0','1','0','0','1','1','1','0'),
            ('1','0','1','1','1','1','0','1','0','1','0','0','0','0'),
            ('1','0','1','1','1','1','0','1','0','1','0','0','1','0'),
            ('1','0','1','1','1','1','0','1','0','1','0','1','0','0'),
            ('1','0','1','1','1','1','0','1','0','1','0','1','1','0'),
            ('1','0','1','1','1','1','0','1','0','1','1','0','0','0'),
            ('1','0','1','1','1','1','0','1','0','1','1','0','1','0'),
            ('1','0','1','1','1','1','0','1','0','1','1','1','0','0'),
            ('1','0','1','1','1','1','0','1','0','1','1','1','1','0'),
            ('1','0','1','1','1','1','0','1','1','0','0','0','0','0'),
            ('1','0','1','1','1','1','0','1','1','0','0','0','1','0'),
            ('1','0','1','1','1','1','0','1','1','0','0','1','0','0'),
            ('1','0','1','1','1','1','0','1','1','0','0','1','1','0'),
            ('1','0','1','1','1','1','0','1','1','0','1','0','0','0'),
            ('1','0','1','1','1','1','0','1','1','0','1','0','1','0'),
            ('1','0','1','1','1','1','0','1','1','0','1','1','0','0'),
            ('1','0','1','1','1','1','0','1','1','0','1','1','1','0'),
            ('1','0','1','1','1','1','0','1','1','1','0','0','0','0'),
            ('1','0','1','1','1','1','0','1','1','1','0','0','1','0'),
            ('1','0','1','1','1','1','0','1','1','1','0','1','0','0'),
            ('1','0','1','1','1','1','0','1','1','1','0','1','1','0'),
            ('1','0','1','1','1','1','0','1','1','1','1','0','0','0'),
            ('1','0','1','1','1','1','0','1','1','1','1','0','1','0'),
            ('1','0','1','1','1','1','0','1','1','1','1','1','0','0'),
            ('1','0','1','1','1','1','0','1','1','1','1','1','1','0'),
            ('1','0','1','1','1','1','1','0','0','0','0','0','0','0'),
            ('1','0','1','1','1','1','1','0','0','0','0','0','1','0'),
            ('1','0','1','1','1','1','1','0','0','0','0','1','0','0'),
            ('1','0','1','1','1','1','1','0','0','0','0','1','1','0'),
            ('1','0','1','1','1','1','1','0','0','0','1','0','0','0'),
            ('1','0','1','1','1','1','1','0','0','0','1','0','1','0'),
            ('1','0','1','1','1','1','1','0','0','0','1','1','0','0'),
            ('1','0','1','1','1','1','1','0','0','0','1','1','1','0'),
            ('1','0','1','1','1','1','1','0','0','1','0','0','0','0'),
            ('1','0','1','1','1','1','1','0','0','1','0','0','1','0'),
            ('1','0','1','1','1','1','1','0','0','1','0','1','0','0'),
            ('1','0','1','1','1','1','1','0','0','1','0','1','1','0'),
            ('1','0','1','1','1','1','1','0','0','1','1','0','0','0'),
            ('1','0','1','1','1','1','1','0','0','1','1','0','1','0'),
            ('1','0','1','1','1','1','1','0','0','1','1','1','0','0'),
            ('1','0','1','1','1','1','1','0','0','1','1','1','1','0'),
            ('1','0','1','1','1','1','1','0','1','0','0','0','0','0'),
            ('1','0','1','1','1','1','1','0','1','0','0','0','1','0'),
            ('1','0','1','1','1','1','1','0','1','0','0','1','0','0'),
            ('1','0','1','1','1','1','1','0','1','0','0','1','1','0'),
            ('1','0','1','1','1','1','1','0','1','0','1','0','0','0'),
            ('1','0','1','1','1','1','1','0','1','0','1','0','1','0'),
            ('1','0','1','1','1','1','1','0','1','0','1','1','0','0'),
            ('1','0','1','1','1','1','1','0','1','0','1','1','1','0'),
            ('1','0','1','1','1','1','1','0','1','1','0','0','0','0'),
            ('1','0','1','1','1','1','1','0','1','1','0','0','1','0'),
            ('1','0','1','1','1','1','1','0','1','1','0','1','0','0'),
            ('1','0','1','1','1','1','1','0','1','1','0','1','1','0'),
            ('1','0','1','1','1','1','1','0','1','1','1','0','0','0'),
            ('1','0','1','1','1','1','1','0','1','1','1','0','1','0'),
            ('1','0','1','1','1','1','1','0','1','1','1','1','0','0'),
            ('1','0','1','1','1','1','1','0','1','1','1','1','1','0'),
            ('1','0','1','1','1','1','1','1','0','0','0','0','0','0'),
            ('1','0','1','1','1','1','1','1','0','0','0','0','1','0'),
            ('1','0','1','1','1','1','1','1','0','0','0','1','0','0'),
            ('1','0','1','1','1','1','1','1','0','0','0','1','1','0'),
            ('1','0','1','1','1','1','1','1','0','0','1','0','0','0'),
            ('1','0','1','1','1','1','1','1','0','0','1','0','1','0'),
            ('1','0','1','1','1','1','1','1','0','0','1','1','0','0'),
            ('1','0','1','1','1','1','1','1','0','0','1','1','1','0'),
            ('1','0','1','1','1','1','1','1','0','1','0','0','0','0'),
            ('1','0','1','1','1','1','1','1','0','1','0','0','1','0'),
            ('1','0','1','1','1','1','1','1','0','1','0','1','0','0'),
            ('1','0','1','1','1','1','1','1','0','1','0','1','1','0'),
            ('1','0','1','1','1','1','1','1','0','1','1','0','0','0'),
            ('1','0','1','1','1','1','1','1','0','1','1','0','1','0'),
            ('1','0','1','1','1','1','1','1','0','1','1','1','0','0'),
            ('1','0','1','1','1','1','1','1','0','1','1','1','1','0'),
            ('1','0','1','1','1','1','1','1','1','0','0','0','0','0'),
            ('1','0','1','1','1','1','1','1','1','0','0','0','1','0'),
            ('1','0','1','1','1','1','1','1','1','0','0','1','0','0'),
            ('1','0','1','1','1','1','1','1','1','0','0','1','1','0'),
            ('1','0','1','1','1','1','1','1','1','0','1','0','0','0'),
            ('1','0','1','1','1','1','1','1','1','0','1','0','1','0'),
            ('1','0','1','1','1','1','1','1','1','0','1','1','0','0'),
            ('1','0','1','1','1','1','1','1','1','0','1','1','1','0'),
            ('1','0','1','1','1','1','1','1','1','1','0','0','0','0'),
            ('1','0','1','1','1','1','1','1','1','1','0','0','1','0'),
            ('1','0','1','1','1','1','1','1','1','1','0','1','0','0'),
            ('1','0','1','1','1','1','1','1','1','1','0','1','1','0'),
            ('1','0','1','1','1','1','1','1','1','1','1','0','0','0'),
            ('1','0','1','1','1','1','1','1','1','1','1','0','1','0'),
            ('1','0','1','1','1','1','1','1','1','1','1','1','0','0'),
            ('1','0','1','1','1','1','1','1','1','1','1','1','1','0'),
            ('1','1','0','0','0','0','0','0','0','0','0','0','0','0'),
            ('1','1','0','0','0','0','0','0','0','0','0','0','1','0'),
            ('1','1','0','0','0','0','0','0','0','0','0','1','0','0'),
            ('1','1','0','0','0','0','0','0','0','0','0','1','1','0'),
            ('1','1','0','0','0','0','0','0','0','0','1','0','0','0'),
            ('1','1','0','0','0','0','0','0','0','0','1','0','1','0'),
            ('1','1','0','0','0','0','0','0','0','0','1','1','0','0'),
            ('1','1','0','0','0','0','0','0','0','0','1','1','1','0'),
            ('1','1','0','0','0','0','0','0','0','1','0','0','0','0'),
            ('1','1','0','0','0','0','0','0','0','1','0','0','1','0'),
            ('1','1','0','0','0','0','0','0','0','1','0','1','0','0'),
            ('1','1','0','0','0','0','0','0','0','1','0','1','1','0'),
            ('1','1','0','0','0','0','0','0','0','1','1','0','0','0'),
            ('1','1','0','0','0','0','0','0','0','1','1','0','1','0'),
            ('1','1','0','0','0','0','0','0','0','1','1','1','0','0'),
            ('1','1','0','0','0','0','0','0','0','1','1','1','1','0'),
            ('1','1','0','0','0','0','0','0','1','0','0','0','0','0'),
            ('1','1','0','0','0','0','0','0','1','0','0','0','1','0'),
            ('1','1','0','0','0','0','0','0','1','0','0','1','0','0'),
            ('1','1','0','0','0','0','0','0','1','0','0','1','1','0'),
            ('1','1','0','0','0','0','0','0','1','0','1','0','0','0'),
            ('1','1','0','0','0','0','0','0','1','0','1','0','1','0'),
            ('1','1','0','0','0','0','0','0','1','0','1','1','0','0'),
            ('1','1','0','0','0','0','0','0','1','0','1','1','1','0'),
            ('1','1','0','0','0','0','0','0','1','1','0','0','0','0'),
            ('1','1','0','0','0','0','0','0','1','1','0','0','1','0'),
            ('1','1','0','0','0','0','0','0','1','1','0','1','0','0'),
            ('1','1','0','0','0','0','0','0','1','1','0','1','1','0'),
            ('1','1','0','0','0','0','0','0','1','1','1','0','0','0'),
            ('1','1','0','0','0','0','0','0','1','1','1','0','1','0'),
            ('1','1','0','0','0','0','0','0','1','1','1','1','0','0'),
            ('1','1','0','0','0','0','0','0','1','1','1','1','1','0'),
            ('1','1','0','0','0','0','0','1','0','0','0','0','0','0'),
            ('1','1','0','0','0','0','0','1','0','0','0','0','1','0'),
            ('1','1','0','0','0','0','0','1','0','0','0','1','0','0'),
            ('1','1','0','0','0','0','0','1','0','0','0','1','1','0'),
            ('1','1','0','0','0','0','0','1','0','0','1','0','0','0'),
            ('1','1','0','0','0','0','0','1','0','0','1','0','1','0'),
            ('1','1','0','0','0','0','0','1','0','0','1','1','0','0'),
            ('1','1','0','0','0','0','0','1','0','0','1','1','1','0'),
            ('1','1','0','0','0','0','0','1','0','1','0','0','0','0'),
            ('1','1','0','0','0','0','0','1','0','1','0','0','1','0'),
            ('1','1','0','0','0','0','0','1','0','1','0','1','0','0'),
            ('1','1','0','0','0','0','0','1','0','1','0','1','1','0'),
            ('1','1','0','0','0','0','0','1','0','1','1','0','0','0'),
            ('1','1','0','0','0','0','0','1','0','1','1','0','1','0'),
            ('1','1','0','0','0','0','0','1','0','1','1','1','0','0'),
            ('1','1','0','0','0','0','0','1','0','1','1','1','1','0'),
            ('1','1','0','0','0','0','0','1','1','0','0','0','0','0'),
            ('1','1','0','0','0','0','0','1','1','0','0','0','1','0'),
            ('1','1','0','0','0','0','0','1','1','0','0','1','0','0'),
            ('1','1','0','0','0','0','0','1','1','0','0','1','1','0'),
            ('1','1','0','0','0','0','0','1','1','0','1','0','0','0'),
            ('1','1','0','0','0','0','0','1','1','0','1','0','1','0'),
            ('1','1','0','0','0','0','0','1','1','0','1','1','0','0'),
            ('1','1','0','0','0','0','0','1','1','0','1','1','1','0'),
            ('1','1','0','0','0','0','0','1','1','1','0','0','0','0'),
            ('1','1','0','0','0','0','0','1','1','1','0','0','1','0'),
            ('1','1','0','0','0','0','0','1','1','1','0','1','0','0'),
            ('1','1','0','0','0','0','0','1','1','1','0','1','1','0'),
            ('1','1','0','0','0','0','0','1','1','1','1','0','0','0'),
            ('1','1','0','0','0','0','0','1','1','1','1','0','1','0'),
            ('1','1','0','0','0','0','0','1','1','1','1','1','0','0'),
            ('1','1','0','0','0','0','0','1','1','1','1','1','1','0'),
            ('1','1','0','0','0','0','1','0','0','0','0','0','0','0'),
            ('1','1','0','0','0','0','1','0','0','0','0','0','1','0'),
            ('1','1','0','0','0','0','1','0','0','0','0','1','0','0'),
            ('1','1','0','0','0','0','1','0','0','0','0','1','1','0'),
            ('1','1','0','0','0','0','1','0','0','0','1','0','0','0'),
            ('1','1','0','0','0','0','1','0','0','0','1','0','1','0'),
            ('1','1','0','0','0','0','1','0','0','0','1','1','0','0'),
            ('1','1','0','0','0','0','1','0','0','0','1','1','1','0'),
            ('1','1','0','0','0','0','1','0','0','1','0','0','0','0'),
            ('1','1','0','0','0','0','1','0','0','1','0','0','1','0'),
            ('1','1','0','0','0','0','1','0','0','1','0','1','0','0'),
            ('1','1','0','0','0','0','1','0','0','1','0','1','1','0'),
            ('1','1','0','0','0','0','1','0','0','1','1','0','0','0'),
            ('1','1','0','0','0','0','1','0','0','1','1','0','1','0'),
            ('1','1','0','0','0','0','1','0','0','1','1','1','0','0'),
            ('1','1','0','0','0','0','1','0','0','1','1','1','1','0'),
            ('1','1','0','0','0','0','1','0','1','0','0','0','0','0'),
            ('1','1','0','0','0','0','1','0','1','0','0','0','1','0'),
            ('1','1','0','0','0','0','1','0','1','0','0','1','0','0'),
            ('1','1','0','0','0','0','1','0','1','0','0','1','1','0'),
            ('1','1','0','0','0','0','1','0','1','0','1','0','0','0'),
            ('1','1','0','0','0','0','1','0','1','0','1','0','1','0'),
            ('1','1','0','0','0','0','1','0','1','0','1','1','0','0'),
            ('1','1','0','0','0','0','1','0','1','0','1','1','1','0'),
            ('1','1','0','0','0','0','1','0','1','1','0','0','0','0'),
            ('1','1','0','0','0','0','1','0','1','1','0','0','1','0'),
            ('1','1','0','0','0','0','1','0','1','1','0','1','0','0'),
            ('1','1','0','0','0','0','1','0','1','1','0','1','1','0'),
            ('1','1','0','0','0','0','1','0','1','1','1','0','0','0'),
            ('1','1','0','0','0','0','1','0','1','1','1','0','1','0'),
            ('1','1','0','0','0','0','1','0','1','1','1','1','0','0'),
            ('1','1','0','0','0','0','1','0','1','1','1','1','1','0'),
            ('1','1','0','0','0','0','1','1','0','0','0','0','0','0'),
            ('1','1','0','0','0','0','1','1','0','0','0','0','1','0'),
            ('1','1','0','0','0','0','1','1','0','0','0','1','0','0'),
            ('1','1','0','0','0','0','1','1','0','0','0','1','1','0'),
            ('1','1','0','0','0','0','1','1','0','0','1','0','0','0'),
            ('1','1','0','0','0','0','1','1','0','0','1','0','1','0'),
            ('1','1','0','0','0','0','1','1','0','0','1','1','0','0'),
            ('1','1','0','0','0','0','1','1','0','0','1','1','1','0'),
            ('1','1','0','0','0','0','1','1','0','1','0','0','0','0'),
            ('1','1','0','0','0','0','1','1','0','1','0','0','1','0'),
            ('1','1','0','0','0','0','1','1','0','1','0','1','0','0'),
            ('1','1','0','0','0','0','1','1','0','1','0','1','1','0'),
            ('1','1','0','0','0','0','1','1','0','1','1','0','0','0'),
            ('1','1','0','0','0','0','1','1','0','1','1','0','1','0'),
            ('1','1','0','0','0','0','1','1','0','1','1','1','0','0'),
            ('1','1','0','0','0','0','1','1','0','1','1','1','1','0'),
            ('1','1','0','0','0','0','1','1','1','0','0','0','0','0'),
            ('1','1','0','0','0','0','1','1','1','0','0','0','1','0'),
            ('1','1','0','0','0','0','1','1','1','0','0','1','0','0'),
            ('1','1','0','0','0','0','1','1','1','0','0','1','1','0'),
            ('1','1','0','0','0','0','1','1','1','0','1','0','0','0'),
            ('1','1','0','0','0','0','1','1','1','0','1','0','1','0'),
            ('1','1','0','0','0','0','1','1','1','0','1','1','0','0'),
            ('1','1','0','0','0','0','1','1','1','0','1','1','1','0'),
            ('1','1','0','0','0','0','1','1','1','1','0','0','0','0'),
            ('1','1','0','0','0','0','1','1','1','1','0','0','1','0'),
            ('1','1','0','0','0','0','1','1','1','1','0','1','0','0'),
            ('1','1','0','0','0','0','1','1','1','1','0','1','1','0'),
            ('1','1','0','0','0','0','1','1','1','1','1','0','0','0'),
            ('1','1','0','0','0','0','1','1','1','1','1','0','1','0'),
            ('1','1','0','0','0','0','1','1','1','1','1','1','0','0'),
            ('1','1','0','0','0','0','1','1','1','1','1','1','1','0'),
            ('1','1','0','0','0','1','0','0','0','0','0','0','0','0'),
            ('1','1','0','0','0','1','0','0','0','0','0','0','1','0'),
            ('1','1','0','0','0','1','0','0','0','0','0','1','0','0'),
            ('1','1','0','0','0','1','0','0','0','0','0','1','1','0'),
            ('1','1','0','0','0','1','0','0','0','0','1','0','0','0'),
            ('1','1','0','0','0','1','0','0','0','0','1','0','1','0'),
            ('1','1','0','0','0','1','0','0','0','0','1','1','0','0'),
            ('1','1','0','0','0','1','0','0','0','0','1','1','1','0'),
            ('1','1','0','0','0','1','0','0','0','1','0','0','0','0'),
            ('1','1','0','0','0','1','0','0','0','1','0','0','1','0'),
            ('1','1','0','0','0','1','0','0','0','1','0','1','0','0'),
            ('1','1','0','0','0','1','0','0','0','1','0','1','1','0'),
            ('1','1','0','0','0','1','0','0','0','1','1','0','0','0'),
            ('1','1','0','0','0','1','0','0','0','1','1','0','1','0'),
            ('1','1','0','0','0','1','0','0','0','1','1','1','0','0'),
            ('1','1','0','0','0','1','0','0','0','1','1','1','1','0'),
            ('1','1','0','0','0','1','0','0','1','0','0','0','0','0'),
            ('1','1','0','0','0','1','0','0','1','0','0','0','1','0'),
            ('1','1','0','0','0','1','0','0','1','0','0','1','0','0'),
            ('1','1','0','0','0','1','0','0','1','0','0','1','1','0'),
            ('1','1','0','0','0','1','0','0','1','0','1','0','0','0'),
            ('1','1','0','0','0','1','0','0','1','0','1','0','1','0'),
            ('1','1','0','0','0','1','0','0','1','0','1','1','0','0'),
            ('1','1','0','0','0','1','0','0','1','0','1','1','1','0'),
            ('1','1','0','0','0','1','0','0','1','1','0','0','0','0'),
            ('1','1','0','0','0','1','0','0','1','1','0','0','1','0'),
            ('1','1','0','0','0','1','0','0','1','1','0','1','0','0'),
            ('1','1','0','0','0','1','0','0','1','1','0','1','1','0'),
            ('1','1','0','0','0','1','0','0','1','1','1','0','0','0'),
            ('1','1','0','0','0','1','0','0','1','1','1','0','1','0'),
            ('1','1','0','0','0','1','0','0','1','1','1','1','0','0'),
            ('1','1','0','0','0','1','0','0','1','1','1','1','1','0'),
            ('1','1','0','0','0','1','0','1','0','0','0','0','0','0'),
            ('1','1','0','0','0','1','0','1','0','0','0','0','1','0'),
            ('1','1','0','0','0','1','0','1','0','0','0','1','0','0'),
            ('1','1','0','0','0','1','0','1','0','0','0','1','1','0'),
            ('1','1','0','0','0','1','0','1','0','0','1','0','0','0'),
            ('1','1','0','0','0','1','0','1','0','0','1','0','1','0'),
            ('1','1','0','0','0','1','0','1','0','0','1','1','0','0'),
            ('1','1','0','0','0','1','0','1','0','0','1','1','1','0'),
            ('1','1','0','0','0','1','0','1','0','1','0','0','0','0'),
            ('1','1','0','0','0','1','0','1','0','1','0','0','1','0'),
            ('1','1','0','0','0','1','0','1','0','1','0','1','0','0'),
            ('1','1','0','0','0','1','0','1','0','1','0','1','1','0'),
            ('1','1','0','0','0','1','0','1','0','1','1','0','0','0'),
            ('1','1','0','0','0','1','0','1','0','1','1','0','1','0'),
            ('1','1','0','0','0','1','0','1','0','1','1','1','0','0'),
            ('1','1','0','0','0','1','0','1','0','1','1','1','1','0'),
            ('1','1','0','0','0','1','0','1','1','0','0','0','0','0'),
            ('1','1','0','0','0','1','0','1','1','0','0','0','1','0'),
            ('1','1','0','0','0','1','0','1','1','0','0','1','0','0'),
            ('1','1','0','0','0','1','0','1','1','0','0','1','1','0'),
            ('1','1','0','0','0','1','0','1','1','0','1','0','0','0'),
            ('1','1','0','0','0','1','0','1','1','0','1','0','1','0'),
            ('1','1','0','0','0','1','0','1','1','0','1','1','0','0'),
            ('1','1','0','0','0','1','0','1','1','0','1','1','1','0'),
            ('1','1','0','0','0','1','0','1','1','1','0','0','0','0'),
            ('1','1','0','0','0','1','0','1','1','1','0','0','1','0'),
            ('1','1','0','0','0','1','0','1','1','1','0','1','0','0'),
            ('1','1','0','0','0','1','0','1','1','1','0','1','1','0'),
            ('1','1','0','0','0','1','0','1','1','1','1','0','0','0'),
            ('1','1','0','0','0','1','0','1','1','1','1','0','1','0'),
            ('1','1','0','0','0','1','0','1','1','1','1','1','0','0'),
            ('1','1','0','0','0','1','0','1','1','1','1','1','1','0'),
            ('1','1','0','0','0','1','1','0','0','0','0','0','0','0'),
            ('1','1','0','0','0','1','1','0','0','0','0','0','1','0'),
            ('1','1','0','0','0','1','1','0','0','0','0','1','0','0'),
            ('1','1','0','0','0','1','1','0','0','0','0','1','1','0'),
            ('1','1','0','0','0','1','1','0','0','0','1','0','0','0'),
            ('1','1','0','0','0','1','1','0','0','0','1','0','1','0'),
            ('1','1','0','0','0','1','1','0','0','0','1','1','0','0'),
            ('1','1','0','0','0','1','1','0','0','0','1','1','1','0'),
            ('1','1','0','0','0','1','1','0','0','1','0','0','0','0'),
            ('1','1','0','0','0','1','1','0','0','1','0','0','1','0'),
            ('1','1','0','0','0','1','1','0','0','1','0','1','0','0'),
            ('1','1','0','0','0','1','1','0','0','1','0','1','1','0'),
            ('1','1','0','0','0','1','1','0','0','1','1','0','0','0'),
            ('1','1','0','0','0','1','1','0','0','1','1','0','1','0'),
            ('1','1','0','0','0','1','1','0','0','1','1','1','0','0'),
            ('1','1','0','0','0','1','1','0','0','1','1','1','1','0'),
            ('1','1','0','0','0','1','1','0','1','0','0','0','0','0'),
            ('1','1','0','0','0','1','1','0','1','0','0','0','1','0'),
            ('1','1','0','0','0','1','1','0','1','0','0','1','0','0'),
            ('1','1','0','0','0','1','1','0','1','0','0','1','1','0'),
            ('1','1','0','0','0','1','1','0','1','0','1','0','0','0'),
            ('1','1','0','0','0','1','1','0','1','0','1','0','1','0'),
            ('1','1','0','0','0','1','1','0','1','0','1','1','0','0'),
            ('1','1','0','0','0','1','1','0','1','0','1','1','1','0'),
            ('1','1','0','0','0','1','1','0','1','1','0','0','0','0'),
            ('1','1','0','0','0','1','1','0','1','1','0','0','1','0'),
            ('1','1','0','0','0','1','1','0','1','1','0','1','0','0'),
            ('1','1','0','0','0','1','1','0','1','1','0','1','1','0'),
            ('1','1','0','0','0','1','1','0','1','1','1','0','0','0'),
            ('1','1','0','0','0','1','1','0','1','1','1','0','1','0'),
            ('1','1','0','0','0','1','1','0','1','1','1','1','0','0'),
            ('1','1','0','0','0','1','1','0','1','1','1','1','1','0'),
            ('1','1','0','0','0','1','1','1','0','0','0','0','0','0'),
            ('1','1','0','0','0','1','1','1','0','0','0','0','1','0'),
            ('1','1','0','0','0','1','1','1','0','0','0','1','0','0'),
            ('1','1','0','0','0','1','1','1','0','0','0','1','1','0'),
            ('1','1','0','0','0','1','1','1','0','0','1','0','0','0'),
            ('1','1','0','0','0','1','1','1','0','0','1','0','1','0'),
            ('1','1','0','0','0','1','1','1','0','0','1','1','0','0'),
            ('1','1','0','0','0','1','1','1','0','0','1','1','1','0'),
            ('1','1','0','0','0','1','1','1','0','1','0','0','0','0'),
            ('1','1','0','0','0','1','1','1','0','1','0','0','1','0'),
            ('1','1','0','0','0','1','1','1','0','1','0','1','0','0'),
            ('1','1','0','0','0','1','1','1','0','1','0','1','1','0'),
            ('1','1','0','0','0','1','1','1','0','1','1','0','0','0'),
            ('1','1','0','0','0','1','1','1','0','1','1','0','1','0'),
            ('1','1','0','0','0','1','1','1','0','1','1','1','0','0'),
            ('1','1','0','0','0','1','1','1','0','1','1','1','1','0'),
            ('1','1','0','0','0','1','1','1','1','0','0','0','0','0'),
            ('1','1','0','0','0','1','1','1','1','0','0','0','1','0'),
            ('1','1','0','0','0','1','1','1','1','0','0','1','0','0'),
            ('1','1','0','0','0','1','1','1','1','0','0','1','1','0'),
            ('1','1','0','0','0','1','1','1','1','0','1','0','0','0'),
            ('1','1','0','0','0','1','1','1','1','0','1','0','1','0'),
            ('1','1','0','0','0','1','1','1','1','0','1','1','0','0'),
            ('1','1','0','0','0','1','1','1','1','0','1','1','1','0'),
            ('1','1','0','0','0','1','1','1','1','1','0','0','0','0'),
            ('1','1','0','0','0','1','1','1','1','1','0','0','1','0'),
            ('1','1','0','0','0','1','1','1','1','1','0','1','0','0'),
            ('1','1','0','0','0','1','1','1','1','1','0','1','1','0'),
            ('1','1','0','0','0','1','1','1','1','1','1','0','0','0'),
            ('1','1','0','0','0','1','1','1','1','1','1','0','1','0'),
            ('1','1','0','0','0','1','1','1','1','1','1','1','0','0'),
            ('1','1','0','0','0','1','1','1','1','1','1','1','1','0'),
            ('1','1','0','0','1','0','0','0','0','0','0','0','0','0'),
            ('1','1','0','0','1','0','0','0','0','0','0','0','1','0'),
            ('1','1','0','0','1','0','0','0','0','0','0','1','0','0'),
            ('1','1','0','0','1','0','0','0','0','0','0','1','1','0'),
            ('1','1','0','0','1','0','0','0','0','0','1','0','0','0'),
            ('1','1','0','0','1','0','0','0','0','0','1','0','1','0'),
            ('1','1','0','0','1','0','0','0','0','0','1','1','0','0'),
            ('1','1','0','0','1','0','0','0','0','0','1','1','1','0'),
            ('1','1','0','0','1','0','0','0','0','1','0','0','0','0'),
            ('1','1','0','0','1','0','0','0','0','1','0','0','1','0'),
            ('1','1','0','0','1','0','0','0','0','1','0','1','0','0'),
            ('1','1','0','0','1','0','0','0','0','1','0','1','1','0'),
            ('1','1','0','0','1','0','0','0','0','1','1','0','0','0'),
            ('1','1','0','0','1','0','0','0','0','1','1','0','1','0'),
            ('1','1','0','0','1','0','0','0','0','1','1','1','0','0'),
            ('1','1','0','0','1','0','0','0','0','1','1','1','1','0'),
            ('1','1','0','0','1','0','0','0','1','0','0','0','0','0'),
            ('1','1','0','0','1','0','0','0','1','0','0','0','1','0'),
            ('1','1','0','0','1','0','0','0','1','0','0','1','0','0'),
            ('1','1','0','0','1','0','0','0','1','0','0','1','1','0'),
            ('1','1','0','0','1','0','0','0','1','0','1','0','0','0'),
            ('1','1','0','0','1','0','0','0','1','0','1','0','1','0'),
            ('1','1','0','0','1','0','0','0','1','0','1','1','0','0'),
            ('1','1','0','0','1','0','0','0','1','0','1','1','1','0'),
            ('1','1','0','0','1','0','0','0','1','1','0','0','0','0'),
            ('1','1','0','0','1','0','0','0','1','1','0','0','1','0'),
            ('1','1','0','0','1','0','0','0','1','1','0','1','0','0'),
            ('1','1','0','0','1','0','0','0','1','1','0','1','1','0'),
            ('1','1','0','0','1','0','0','0','1','1','1','0','0','0'),
            ('1','1','0','0','1','0','0','0','1','1','1','0','1','0'),
            ('1','1','0','0','1','0','0','0','1','1','1','1','0','0'),
            ('1','1','0','0','1','0','0','0','1','1','1','1','1','0'),
            ('1','1','0','0','1','0','0','1','0','0','0','0','0','0'),
            ('1','1','0','0','1','0','0','1','0','0','0','0','1','0'),
            ('1','1','0','0','1','0','0','1','0','0','0','1','0','0'),
            ('1','1','0','0','1','0','0','1','0','0','0','1','1','0'),
            ('1','1','0','0','1','0','0','1','0','0','1','0','0','0'),
            ('1','1','0','0','1','0','0','1','0','0','1','0','1','0'),
            ('1','1','0','0','1','0','0','1','0','0','1','1','0','0'),
            ('1','1','0','0','1','0','0','1','0','0','1','1','1','0'),
            ('1','1','0','0','1','0','0','1','0','1','0','0','0','0'),
            ('1','1','0','0','1','0','0','1','0','1','0','0','1','0'),
            ('1','1','0','0','1','0','0','1','0','1','0','1','0','0'),
            ('1','1','0','0','1','0','0','1','0','1','0','1','1','0'),
            ('1','1','0','0','1','0','0','1','0','1','1','0','0','0'),
            ('1','1','0','0','1','0','0','1','0','1','1','0','1','0'),
            ('1','1','0','0','1','0','0','1','0','1','1','1','0','0'),
            ('1','1','0','0','1','0','0','1','0','1','1','1','1','0'),
            ('1','1','0','0','1','0','0','1','1','0','0','0','0','0'),
            ('1','1','0','0','1','0','0','1','1','0','0','0','1','0'),
            ('1','1','0','0','1','0','0','1','1','0','0','1','0','0'),
            ('1','1','0','0','1','0','0','1','1','0','0','1','1','0'),
            ('1','1','0','0','1','0','0','1','1','0','1','0','0','0'),
            ('1','1','0','0','1','0','0','1','1','0','1','0','1','0'),
            ('1','1','0','0','1','0','0','1','1','0','1','1','0','0'),
            ('1','1','0','0','1','0','0','1','1','0','1','1','1','0'),
            ('1','1','0','0','1','0','0','1','1','1','0','0','0','0'),
            ('1','1','0','0','1','0','0','1','1','1','0','0','1','0'),
            ('1','1','0','0','1','0','0','1','1','1','0','1','0','0'),
            ('1','1','0','0','1','0','0','1','1','1','0','1','1','0'),
            ('1','1','0','0','1','0','0','1','1','1','1','0','0','0'),
            ('1','1','0','0','1','0','0','1','1','1','1','0','1','0'),
            ('1','1','0','0','1','0','0','1','1','1','1','1','0','0'),
            ('1','1','0','0','1','0','0','1','1','1','1','1','1','0'),
            ('1','1','0','0','1','0','1','0','0','0','0','0','0','0'),
            ('1','1','0','0','1','0','1','0','0','0','0','0','1','0'),
            ('1','1','0','0','1','0','1','0','0','0','0','1','0','0'),
            ('1','1','0','0','1','0','1','0','0','0','0','1','1','0'),
            ('1','1','0','0','1','0','1','0','0','0','1','0','0','0'),
            ('1','1','0','0','1','0','1','0','0','0','1','0','1','0'),
            ('1','1','0','0','1','0','1','0','0','0','1','1','0','0'),
            ('1','1','0','0','1','0','1','0','0','0','1','1','1','0'),
            ('1','1','0','0','1','0','1','0','0','1','0','0','0','0'),
            ('1','1','0','0','1','0','1','0','0','1','0','0','1','0'),
            ('1','1','0','0','1','0','1','0','0','1','0','1','0','0'),
            ('1','1','0','0','1','0','1','0','0','1','0','1','1','0'),
            ('1','1','0','0','1','0','1','0','0','1','1','0','0','0'),
            ('1','1','0','0','1','0','1','0','0','1','1','0','1','0'),
            ('1','1','0','0','1','0','1','0','0','1','1','1','0','0'),
            ('1','1','0','0','1','0','1','0','0','1','1','1','1','0'),
            ('1','1','0','0','1','0','1','0','1','0','0','0','0','0'),
            ('1','1','0','0','1','0','1','0','1','0','0','0','1','0'),
            ('1','1','0','0','1','0','1','0','1','0','0','1','0','0'),
            ('1','1','0','0','1','0','1','0','1','0','0','1','1','0'),
            ('1','1','0','0','1','0','1','0','1','0','1','0','0','0'),
            ('1','1','0','0','1','0','1','0','1','0','1','0','1','0'),
            ('1','1','0','0','1','0','1','0','1','0','1','1','0','0'),
            ('1','1','0','0','1','0','1','0','1','0','1','1','1','0'),
            ('1','1','0','0','1','0','1','0','1','1','0','0','0','0'),
            ('1','1','0','0','1','0','1','0','1','1','0','0','1','0'),
            ('1','1','0','0','1','0','1','0','1','1','0','1','0','0'),
            ('1','1','0','0','1','0','1','0','1','1','0','1','1','0'),
            ('1','1','0','0','1','0','1','0','1','1','1','0','0','0'),
            ('1','1','0','0','1','0','1','0','1','1','1','0','1','0'),
            ('1','1','0','0','1','0','1','0','1','1','1','1','0','0'),
            ('1','1','0','0','1','0','1','0','1','1','1','1','1','0'),
            ('1','1','0','0','1','0','1','1','0','0','0','0','0','0'),
            ('1','1','0','0','1','0','1','1','0','0','0','0','1','0'),
            ('1','1','0','0','1','0','1','1','0','0','0','1','0','0'),
            ('1','1','0','0','1','0','1','1','0','0','0','1','1','0'),
            ('1','1','0','0','1','0','1','1','0','0','1','0','0','0'),
            ('1','1','0','0','1','0','1','1','0','0','1','0','1','0'),
            ('1','1','0','0','1','0','1','1','0','0','1','1','0','0'),
            ('1','1','0','0','1','0','1','1','0','0','1','1','1','0'),
            ('1','1','0','0','1','0','1','1','0','1','0','0','0','0'),
            ('1','1','0','0','1','0','1','1','0','1','0','0','1','0'),
            ('1','1','0','0','1','0','1','1','0','1','0','1','0','0'),
            ('1','1','0','0','1','0','1','1','0','1','0','1','1','0'),
            ('1','1','0','0','1','0','1','1','0','1','1','0','0','0'),
            ('1','1','0','0','1','0','1','1','0','1','1','0','1','0'),
            ('1','1','0','0','1','0','1','1','0','1','1','1','0','0'),
            ('1','1','0','0','1','0','1','1','0','1','1','1','1','0'),
            ('1','1','0','0','1','0','1','1','1','0','0','0','0','0'),
            ('1','1','0','0','1','0','1','1','1','0','0','0','1','0'),
            ('1','1','0','0','1','0','1','1','1','0','0','1','0','0'),
            ('1','1','0','0','1','0','1','1','1','0','0','1','1','0'),
            ('1','1','0','0','1','0','1','1','1','0','1','0','0','0'),
            ('1','1','0','0','1','0','1','1','1','0','1','0','1','0'),
            ('1','1','0','0','1','0','1','1','1','0','1','1','0','0'),
            ('1','1','0','0','1','0','1','1','1','0','1','1','1','0'),
            ('1','1','0','0','1','0','1','1','1','1','0','0','0','0'),
            ('1','1','0','0','1','0','1','1','1','1','0','0','1','0'),
            ('1','1','0','0','1','0','1','1','1','1','0','1','0','0'),
            ('1','1','0','0','1','0','1','1','1','1','0','1','1','0'),
            ('1','1','0','0','1','0','1','1','1','1','1','0','0','0'),
            ('1','1','0','0','1','0','1','1','1','1','1','0','1','0'),
            ('1','1','0','0','1','0','1','1','1','1','1','1','0','0'),
            ('1','1','0','0','1','0','1','1','1','1','1','1','1','0'),
            ('1','1','0','0','1','1','0','0','0','0','0','0','0','0'),
            ('1','1','0','0','1','1','0','0','0','0','0','0','1','0'),
            ('1','1','0','0','1','1','0','0','0','0','0','1','0','0'),
            ('1','1','0','0','1','1','0','0','0','0','0','1','1','0'),
            ('1','1','0','0','1','1','0','0','0','0','1','0','0','0'),
            ('1','1','0','0','1','1','0','0','0','0','1','0','1','0'),
            ('1','1','0','0','1','1','0','0','0','0','1','1','0','0'),
            ('1','1','0','0','1','1','0','0','0','0','1','1','1','0'),
            ('1','1','0','0','1','1','0','0','0','1','0','0','0','0'),
            ('1','1','0','0','1','1','0','0','0','1','0','0','1','0'),
            ('1','1','0','0','1','1','0','0','0','1','0','1','0','0'),
            ('1','1','0','0','1','1','0','0','0','1','0','1','1','0'),
            ('1','1','0','0','1','1','0','0','0','1','1','0','0','0'),
            ('1','1','0','0','1','1','0','0','0','1','1','0','1','0'),
            ('1','1','0','0','1','1','0','0','0','1','1','1','0','0'),
            ('1','1','0','0','1','1','0','0','0','1','1','1','1','0'),
            ('1','1','0','0','1','1','0','0','1','0','0','0','0','0'),
            ('1','1','0','0','1','1','0','0','1','0','0','0','1','0'),
            ('1','1','0','0','1','1','0','0','1','0','0','1','0','0'),
            ('1','1','0','0','1','1','0','0','1','0','0','1','1','0'),
            ('1','1','0','0','1','1','0','0','1','0','1','0','0','0'),
            ('1','1','0','0','1','1','0','0','1','0','1','0','1','0'),
            ('1','1','0','0','1','1','0','0','1','0','1','1','0','0'),
            ('1','1','0','0','1','1','0','0','1','0','1','1','1','0'),
            ('1','1','0','0','1','1','0','0','1','1','0','0','0','0'),
            ('1','1','0','0','1','1','0','0','1','1','0','0','1','0'),
            ('1','1','0','0','1','1','0','0','1','1','0','1','0','0'),
            ('1','1','0','0','1','1','0','0','1','1','0','1','1','0'),
            ('1','1','0','0','1','1','0','0','1','1','1','0','0','0'),
            ('1','1','0','0','1','1','0','0','1','1','1','0','1','0'),
            ('1','1','0','0','1','1','0','0','1','1','1','1','0','0'),
            ('1','1','0','0','1','1','0','0','1','1','1','1','1','0'),
            ('1','1','0','0','1','1','0','1','0','0','0','0','0','0'),
            ('1','1','0','0','1','1','0','1','0','0','0','0','1','0'),
            ('1','1','0','0','1','1','0','1','0','0','0','1','0','0'),
            ('1','1','0','0','1','1','0','1','0','0','0','1','1','0'),
            ('1','1','0','0','1','1','0','1','0','0','1','0','0','0'),
            ('1','1','0','0','1','1','0','1','0','0','1','0','1','0'),
            ('1','1','0','0','1','1','0','1','0','0','1','1','0','0'),
            ('1','1','0','0','1','1','0','1','0','0','1','1','1','0'),
            ('1','1','0','0','1','1','0','1','0','1','0','0','0','0'),
            ('1','1','0','0','1','1','0','1','0','1','0','0','1','0'),
            ('1','1','0','0','1','1','0','1','0','1','0','1','0','0'),
            ('1','1','0','0','1','1','0','1','0','1','0','1','1','0'),
            ('1','1','0','0','1','1','0','1','0','1','1','0','0','0'),
            ('1','1','0','0','1','1','0','1','0','1','1','0','1','0'),
            ('1','1','0','0','1','1','0','1','0','1','1','1','0','0'),
            ('1','1','0','0','1','1','0','1','0','1','1','1','1','0'),
            ('1','1','0','0','1','1','0','1','1','0','0','0','0','0'),
            ('1','1','0','0','1','1','0','1','1','0','0','0','1','0'),
            ('1','1','0','0','1','1','0','1','1','0','0','1','0','0'),
            ('1','1','0','0','1','1','0','1','1','0','0','1','1','0'),
            ('1','1','0','0','1','1','0','1','1','0','1','0','0','0'),
            ('1','1','0','0','1','1','0','1','1','0','1','0','1','0'),
            ('1','1','0','0','1','1','0','1','1','0','1','1','0','0'),
            ('1','1','0','0','1','1','0','1','1','0','1','1','1','0'),
            ('1','1','0','0','1','1','0','1','1','1','0','0','0','0'),
            ('1','1','0','0','1','1','0','1','1','1','0','0','1','0'),
            ('1','1','0','0','1','1','0','1','1','1','0','1','0','0'),
            ('1','1','0','0','1','1','0','1','1','1','0','1','1','0'),
            ('1','1','0','0','1','1','0','1','1','1','1','0','0','0'),
            ('1','1','0','0','1','1','0','1','1','1','1','0','1','0'),
            ('1','1','0','0','1','1','0','1','1','1','1','1','0','0'),
            ('1','1','0','0','1','1','0','1','1','1','1','1','1','0'),
            ('1','1','0','0','1','1','1','0','0','0','0','0','0','0'),
            ('1','1','0','0','1','1','1','0','0','0','0','0','1','0'),
            ('1','1','0','0','1','1','1','0','0','0','0','1','0','0'),
            ('1','1','0','0','1','1','1','0','0','0','0','1','1','0'),
            ('1','1','0','0','1','1','1','0','0','0','1','0','0','0'),
            ('1','1','0','0','1','1','1','0','0','0','1','0','1','0'),
            ('1','1','0','0','1','1','1','0','0','0','1','1','0','0'),
            ('1','1','0','0','1','1','1','0','0','0','1','1','1','0'),
            ('1','1','0','0','1','1','1','0','0','1','0','0','0','0'),
            ('1','1','0','0','1','1','1','0','0','1','0','0','1','0'),
            ('1','1','0','0','1','1','1','0','0','1','0','1','0','0'),
            ('1','1','0','0','1','1','1','0','0','1','0','1','1','0'),
            ('1','1','0','0','1','1','1','0','0','1','1','0','0','0'),
            ('1','1','0','0','1','1','1','0','0','1','1','0','1','0'),
            ('1','1','0','0','1','1','1','0','0','1','1','1','0','0'),
            ('1','1','0','0','1','1','1','0','0','1','1','1','1','0'),
            ('1','1','0','0','1','1','1','0','1','0','0','0','0','0'),
            ('1','1','0','0','1','1','1','0','1','0','0','0','1','0'),
            ('1','1','0','0','1','1','1','0','1','0','0','1','0','0'),
            ('1','1','0','0','1','1','1','0','1','0','0','1','1','0'),
            ('1','1','0','0','1','1','1','0','1','0','1','0','0','0'),
            ('1','1','0','0','1','1','1','0','1','0','1','0','1','0'),
            ('1','1','0','0','1','1','1','0','1','0','1','1','0','0'),
            ('1','1','0','0','1','1','1','0','1','0','1','1','1','0'),
            ('1','1','0','0','1','1','1','0','1','1','0','0','0','0'),
            ('1','1','0','0','1','1','1','0','1','1','0','0','1','0'),
            ('1','1','0','0','1','1','1','0','1','1','0','1','0','0'),
            ('1','1','0','0','1','1','1','0','1','1','0','1','1','0'),
            ('1','1','0','0','1','1','1','0','1','1','1','0','0','0'),
            ('1','1','0','0','1','1','1','0','1','1','1','0','1','0'),
            ('1','1','0','0','1','1','1','0','1','1','1','1','0','0'),
            ('1','1','0','0','1','1','1','0','1','1','1','1','1','0'),
            ('1','1','0','0','1','1','1','1','0','0','0','0','0','0'),
            ('1','1','0','0','1','1','1','1','0','0','0','0','1','0'),
            ('1','1','0','0','1','1','1','1','0','0','0','1','0','0'),
            ('1','1','0','0','1','1','1','1','0','0','0','1','1','0'),
            ('1','1','0','0','1','1','1','1','0','0','1','0','0','0'),
            ('1','1','0','0','1','1','1','1','0','0','1','0','1','0'),
            ('1','1','0','0','1','1','1','1','0','0','1','1','0','0'),
            ('1','1','0','0','1','1','1','1','0','0','1','1','1','0'),
            ('1','1','0','0','1','1','1','1','0','1','0','0','0','0'),
            ('1','1','0','0','1','1','1','1','0','1','0','0','1','0'),
            ('1','1','0','0','1','1','1','1','0','1','0','1','0','0'),
            ('1','1','0','0','1','1','1','1','0','1','0','1','1','0'),
            ('1','1','0','0','1','1','1','1','0','1','1','0','0','0'),
            ('1','1','0','0','1','1','1','1','0','1','1','0','1','0'),
            ('1','1','0','0','1','1','1','1','0','1','1','1','0','0'),
            ('1','1','0','0','1','1','1','1','0','1','1','1','1','0'),
            ('1','1','0','0','1','1','1','1','1','0','0','0','0','0'),
            ('1','1','0','0','1','1','1','1','1','0','0','0','1','0'),
            ('1','1','0','0','1','1','1','1','1','0','0','1','0','0'),
            ('1','1','0','0','1','1','1','1','1','0','0','1','1','0'),
            ('1','1','0','0','1','1','1','1','1','0','1','0','0','0'),
            ('1','1','0','0','1','1','1','1','1','0','1','0','1','0'),
            ('1','1','0','0','1','1','1','1','1','0','1','1','0','0'),
            ('1','1','0','0','1','1','1','1','1','0','1','1','1','0'),
            ('1','1','0','0','1','1','1','1','1','1','0','0','0','0'),
            ('1','1','0','0','1','1','1','1','1','1','0','0','1','0'),
            ('1','1','0','0','1','1','1','1','1','1','0','1','0','0'),
            ('1','1','0','0','1','1','1','1','1','1','0','1','1','0'),
            ('1','1','0','0','1','1','1','1','1','1','1','0','0','0'),
            ('1','1','0','0','1','1','1','1','1','1','1','0','1','0'),
            ('1','1','0','0','1','1','1','1','1','1','1','1','0','0'),
            ('1','1','0','0','1','1','1','1','1','1','1','1','1','0'),
            ('1','1','0','1','0','0','0','0','0','0','0','0','0','0'),
            ('1','1','0','1','0','0','0','0','0','0','0','0','1','0'),
            ('1','1','0','1','0','0','0','0','0','0','0','1','0','0'),
            ('1','1','0','1','0','0','0','0','0','0','0','1','1','0'),
            ('1','1','0','1','0','0','0','0','0','0','1','0','0','0'),
            ('1','1','0','1','0','0','0','0','0','0','1','0','1','0'),
            ('1','1','0','1','0','0','0','0','0','0','1','1','0','0'),
            ('1','1','0','1','0','0','0','0','0','0','1','1','1','0'),
            ('1','1','0','1','0','0','0','0','0','1','0','0','0','0'),
            ('1','1','0','1','0','0','0','0','0','1','0','0','1','0'),
            ('1','1','0','1','0','0','0','0','0','1','0','1','0','0'),
            ('1','1','0','1','0','0','0','0','0','1','0','1','1','0'),
            ('1','1','0','1','0','0','0','0','0','1','1','0','0','0'),
            ('1','1','0','1','0','0','0','0','0','1','1','0','1','0'),
            ('1','1','0','1','0','0','0','0','0','1','1','1','0','0'),
            ('1','1','0','1','0','0','0','0','0','1','1','1','1','0'),
            ('1','1','0','1','0','0','0','0','1','0','0','0','0','0'),
            ('1','1','0','1','0','0','0','0','1','0','0','0','1','0'),
            ('1','1','0','1','0','0','0','0','1','0','0','1','0','0'),
            ('1','1','0','1','0','0','0','0','1','0','0','1','1','0'),
            ('1','1','0','1','0','0','0','0','1','0','1','0','0','0'),
            ('1','1','0','1','0','0','0','0','1','0','1','0','1','0'),
            ('1','1','0','1','0','0','0','0','1','0','1','1','0','0'),
            ('1','1','0','1','0','0','0','0','1','0','1','1','1','0'),
            ('1','1','0','1','0','0','0','0','1','1','0','0','0','0'),
            ('1','1','0','1','0','0','0','0','1','1','0','0','1','0'),
            ('1','1','0','1','0','0','0','0','1','1','0','1','0','0'),
            ('1','1','0','1','0','0','0','0','1','1','0','1','1','0'),
            ('1','1','0','1','0','0','0','0','1','1','1','0','0','0'),
            ('1','1','0','1','0','0','0','0','1','1','1','0','1','0'),
            ('1','1','0','1','0','0','0','0','1','1','1','1','0','0'),
            ('1','1','0','1','0','0','0','0','1','1','1','1','1','0'),
            ('1','1','0','1','0','0','0','1','0','0','0','0','0','0'),
            ('1','1','0','1','0','0','0','1','0','0','0','0','1','0'),
            ('1','1','0','1','0','0','0','1','0','0','0','1','0','0'),
            ('1','1','0','1','0','0','0','1','0','0','0','1','1','0'),
            ('1','1','0','1','0','0','0','1','0','0','1','0','0','0'),
            ('1','1','0','1','0','0','0','1','0','0','1','0','1','0'),
            ('1','1','0','1','0','0','0','1','0','0','1','1','0','0'),
            ('1','1','0','1','0','0','0','1','0','0','1','1','1','0'),
            ('1','1','0','1','0','0','0','1','0','1','0','0','0','0'),
            ('1','1','0','1','0','0','0','1','0','1','0','0','1','0'),
            ('1','1','0','1','0','0','0','1','0','1','0','1','0','0'),
            ('1','1','0','1','0','0','0','1','0','1','0','1','1','0'),
            ('1','1','0','1','0','0','0','1','0','1','1','0','0','0'),
            ('1','1','0','1','0','0','0','1','0','1','1','0','1','0'),
            ('1','1','0','1','0','0','0','1','0','1','1','1','0','0'),
            ('1','1','0','1','0','0','0','1','0','1','1','1','1','0'),
            ('1','1','0','1','0','0','0','1','1','0','0','0','0','0'),
            ('1','1','0','1','0','0','0','1','1','0','0','0','1','0'),
            ('1','1','0','1','0','0','0','1','1','0','0','1','0','0'),
            ('1','1','0','1','0','0','0','1','1','0','0','1','1','0'),
            ('1','1','0','1','0','0','0','1','1','0','1','0','0','0'),
            ('1','1','0','1','0','0','0','1','1','0','1','0','1','0'),
            ('1','1','0','1','0','0','0','1','1','0','1','1','0','0'),
            ('1','1','0','1','0','0','0','1','1','0','1','1','1','0'),
            ('1','1','0','1','0','0','0','1','1','1','0','0','0','0'),
            ('1','1','0','1','0','0','0','1','1','1','0','0','1','0'),
            ('1','1','0','1','0','0','0','1','1','1','0','1','0','0'),
            ('1','1','0','1','0','0','0','1','1','1','0','1','1','0'),
            ('1','1','0','1','0','0','0','1','1','1','1','0','0','0'),
            ('1','1','0','1','0','0','0','1','1','1','1','0','1','0'),
            ('1','1','0','1','0','0','0','1','1','1','1','1','0','0'),
            ('1','1','0','1','0','0','0','1','1','1','1','1','1','0'),
            ('1','1','0','1','0','0','1','0','0','0','0','0','0','0'),
            ('1','1','0','1','0','0','1','0','0','0','0','0','1','0'),
            ('1','1','0','1','0','0','1','0','0','0','0','1','0','0'),
            ('1','1','0','1','0','0','1','0','0','0','0','1','1','0'),
            ('1','1','0','1','0','0','1','0','0','0','1','0','0','0'),
            ('1','1','0','1','0','0','1','0','0','0','1','0','1','0'),
            ('1','1','0','1','0','0','1','0','0','0','1','1','0','0'),
            ('1','1','0','1','0','0','1','0','0','0','1','1','1','0'),
            ('1','1','0','1','0','0','1','0','0','1','0','0','0','0'),
            ('1','1','0','1','0','0','1','0','0','1','0','0','1','0'),
            ('1','1','0','1','0','0','1','0','0','1','0','1','0','0'),
            ('1','1','0','1','0','0','1','0','0','1','0','1','1','0'),
            ('1','1','0','1','0','0','1','0','0','1','1','0','0','0'),
            ('1','1','0','1','0','0','1','0','0','1','1','0','1','0'),
            ('1','1','0','1','0','0','1','0','0','1','1','1','0','0'),
            ('1','1','0','1','0','0','1','0','0','1','1','1','1','0'),
            ('1','1','0','1','0','0','1','0','1','0','0','0','0','0'),
            ('1','1','0','1','0','0','1','0','1','0','0','0','1','0'),
            ('1','1','0','1','0','0','1','0','1','0','0','1','0','0'),
            ('1','1','0','1','0','0','1','0','1','0','0','1','1','0'),
            ('1','1','0','1','0','0','1','0','1','0','1','0','0','0'),
            ('1','1','0','1','0','0','1','0','1','0','1','0','1','0'),
            ('1','1','0','1','0','0','1','0','1','0','1','1','0','0'),
            ('1','1','0','1','0','0','1','0','1','0','1','1','1','0'),
            ('1','1','0','1','0','0','1','0','1','1','0','0','0','0'),
            ('1','1','0','1','0','0','1','0','1','1','0','0','1','0'),
            ('1','1','0','1','0','0','1','0','1','1','0','1','0','0'),
            ('1','1','0','1','0','0','1','0','1','1','0','1','1','0'),
            ('1','1','0','1','0','0','1','0','1','1','1','0','0','0'),
            ('1','1','0','1','0','0','1','0','1','1','1','0','1','0'),
            ('1','1','0','1','0','0','1','0','1','1','1','1','0','0'),
            ('1','1','0','1','0','0','1','0','1','1','1','1','1','0'),
            ('1','1','0','1','0','0','1','1','0','0','0','0','0','0'),
            ('1','1','0','1','0','0','1','1','0','0','0','0','1','0'),
            ('1','1','0','1','0','0','1','1','0','0','0','1','0','0'),
            ('1','1','0','1','0','0','1','1','0','0','0','1','1','0'),
            ('1','1','0','1','0','0','1','1','0','0','1','0','0','0'),
            ('1','1','0','1','0','0','1','1','0','0','1','0','1','0'),
            ('1','1','0','1','0','0','1','1','0','0','1','1','0','0'),
            ('1','1','0','1','0','0','1','1','0','0','1','1','1','0'),
            ('1','1','0','1','0','0','1','1','0','1','0','0','0','0'),
            ('1','1','0','1','0','0','1','1','0','1','0','0','1','0'),
            ('1','1','0','1','0','0','1','1','0','1','0','1','0','0'),
            ('1','1','0','1','0','0','1','1','0','1','0','1','1','0'),
            ('1','1','0','1','0','0','1','1','0','1','1','0','0','0'),
            ('1','1','0','1','0','0','1','1','0','1','1','0','1','0'),
            ('1','1','0','1','0','0','1','1','0','1','1','1','0','0'),
            ('1','1','0','1','0','0','1','1','0','1','1','1','1','0'),
            ('1','1','0','1','0','0','1','1','1','0','0','0','0','0'),
            ('1','1','0','1','0','0','1','1','1','0','0','0','1','0'),
            ('1','1','0','1','0','0','1','1','1','0','0','1','0','0'),
            ('1','1','0','1','0','0','1','1','1','0','0','1','1','0'),
            ('1','1','0','1','0','0','1','1','1','0','1','0','0','0'),
            ('1','1','0','1','0','0','1','1','1','0','1','0','1','0'),
            ('1','1','0','1','0','0','1','1','1','0','1','1','0','0'),
            ('1','1','0','1','0','0','1','1','1','0','1','1','1','0'),
            ('1','1','0','1','0','0','1','1','1','1','0','0','0','0'),
            ('1','1','0','1','0','0','1','1','1','1','0','0','1','0'),
            ('1','1','0','1','0','0','1','1','1','1','0','1','0','0'),
            ('1','1','0','1','0','0','1','1','1','1','0','1','1','0'),
            ('1','1','0','1','0','0','1','1','1','1','1','0','0','0'),
            ('1','1','0','1','0','0','1','1','1','1','1','0','1','0'),
            ('1','1','0','1','0','0','1','1','1','1','1','1','0','0'),
            ('1','1','0','1','0','0','1','1','1','1','1','1','1','0'),
            ('1','1','0','1','0','1','0','0','0','0','0','0','0','0'),
            ('1','1','0','1','0','1','0','0','0','0','0','0','1','0'),
            ('1','1','0','1','0','1','0','0','0','0','0','1','0','0'),
            ('1','1','0','1','0','1','0','0','0','0','0','1','1','0'),
            ('1','1','0','1','0','1','0','0','0','0','1','0','0','0'),
            ('1','1','0','1','0','1','0','0','0','0','1','0','1','0'),
            ('1','1','0','1','0','1','0','0','0','0','1','1','0','0'),
            ('1','1','0','1','0','1','0','0','0','0','1','1','1','0'),
            ('1','1','0','1','0','1','0','0','0','1','0','0','0','0'),
            ('1','1','0','1','0','1','0','0','0','1','0','0','1','0'),
            ('1','1','0','1','0','1','0','0','0','1','0','1','0','0'),
            ('1','1','0','1','0','1','0','0','0','1','0','1','1','0'),
            ('1','1','0','1','0','1','0','0','0','1','1','0','0','0'),
            ('1','1','0','1','0','1','0','0','0','1','1','0','1','0'),
            ('1','1','0','1','0','1','0','0','0','1','1','1','0','0'),
            ('1','1','0','1','0','1','0','0','0','1','1','1','1','0'),
            ('1','1','0','1','0','1','0','0','1','0','0','0','0','0'),
            ('1','1','0','1','0','1','0','0','1','0','0','0','1','0'),
            ('1','1','0','1','0','1','0','0','1','0','0','1','0','0'),
            ('1','1','0','1','0','1','0','0','1','0','0','1','1','0'),
            ('1','1','0','1','0','1','0','0','1','0','1','0','0','0'),
            ('1','1','0','1','0','1','0','0','1','0','1','0','1','0'),
            ('1','1','0','1','0','1','0','0','1','0','1','1','0','0'),
            ('1','1','0','1','0','1','0','0','1','0','1','1','1','0'),
            ('1','1','0','1','0','1','0','0','1','1','0','0','0','0'),
            ('1','1','0','1','0','1','0','0','1','1','0','0','1','0'),
            ('1','1','0','1','0','1','0','0','1','1','0','1','0','0'),
            ('1','1','0','1','0','1','0','0','1','1','0','1','1','0'),
            ('1','1','0','1','0','1','0','0','1','1','1','0','0','0'),
            ('1','1','0','1','0','1','0','0','1','1','1','0','1','0'),
            ('1','1','0','1','0','1','0','0','1','1','1','1','0','0'),
            ('1','1','0','1','0','1','0','0','1','1','1','1','1','0'),
            ('1','1','0','1','0','1','0','1','0','0','0','0','0','0'),
            ('1','1','0','1','0','1','0','1','0','0','0','0','1','0'),
            ('1','1','0','1','0','1','0','1','0','0','0','1','0','0'),
            ('1','1','0','1','0','1','0','1','0','0','0','1','1','0'),
            ('1','1','0','1','0','1','0','1','0','0','1','0','0','0'),
            ('1','1','0','1','0','1','0','1','0','0','1','0','1','0'),
            ('1','1','0','1','0','1','0','1','0','0','1','1','0','0'),
            ('1','1','0','1','0','1','0','1','0','0','1','1','1','0'),
            ('1','1','0','1','0','1','0','1','0','1','0','0','0','0'),
            ('1','1','0','1','0','1','0','1','0','1','0','0','1','0'),
            ('1','1','0','1','0','1','0','1','0','1','0','1','0','0'),
            ('1','1','0','1','0','1','0','1','0','1','0','1','1','0'),
            ('1','1','0','1','0','1','0','1','0','1','1','0','0','0'),
            ('1','1','0','1','0','1','0','1','0','1','1','0','1','0'),
            ('1','1','0','1','0','1','0','1','0','1','1','1','0','0'),
            ('1','1','0','1','0','1','0','1','0','1','1','1','1','0'),
            ('1','1','0','1','0','1','0','1','1','0','0','0','0','0'),
            ('1','1','0','1','0','1','0','1','1','0','0','0','1','0'),
            ('1','1','0','1','0','1','0','1','1','0','0','1','0','0'),
            ('1','1','0','1','0','1','0','1','1','0','0','1','1','0'),
            ('1','1','0','1','0','1','0','1','1','0','1','0','0','0'),
            ('1','1','0','1','0','1','0','1','1','0','1','0','1','0'),
            ('1','1','0','1','0','1','0','1','1','0','1','1','0','0'),
            ('1','1','0','1','0','1','0','1','1','0','1','1','1','0'),
            ('1','1','0','1','0','1','0','1','1','1','0','0','0','0'),
            ('1','1','0','1','0','1','0','1','1','1','0','0','1','0'),
            ('1','1','0','1','0','1','0','1','1','1','0','1','0','0'),
            ('1','1','0','1','0','1','0','1','1','1','0','1','1','0'),
            ('1','1','0','1','0','1','0','1','1','1','1','0','0','0'),
            ('1','1','0','1','0','1','0','1','1','1','1','0','1','0'),
            ('1','1','0','1','0','1','0','1','1','1','1','1','0','0'),
            ('1','1','0','1','0','1','0','1','1','1','1','1','1','0'),
            ('1','1','0','1','0','1','1','0','0','0','0','0','0','0'),
            ('1','1','0','1','0','1','1','0','0','0','0','0','1','0'),
            ('1','1','0','1','0','1','1','0','0','0','0','1','0','0'),
            ('1','1','0','1','0','1','1','0','0','0','0','1','1','0'),
            ('1','1','0','1','0','1','1','0','0','0','1','0','0','0'),
            ('1','1','0','1','0','1','1','0','0','0','1','0','1','0'),
            ('1','1','0','1','0','1','1','0','0','0','1','1','0','0'),
            ('1','1','0','1','0','1','1','0','0','0','1','1','1','0'),
            ('1','1','0','1','0','1','1','0','0','1','0','0','0','0'),
            ('1','1','0','1','0','1','1','0','0','1','0','0','1','0'),
            ('1','1','0','1','0','1','1','0','0','1','0','1','0','0'),
            ('1','1','0','1','0','1','1','0','0','1','0','1','1','0'),
            ('1','1','0','1','0','1','1','0','0','1','1','0','0','0'),
            ('1','1','0','1','0','1','1','0','0','1','1','0','1','0'),
            ('1','1','0','1','0','1','1','0','0','1','1','1','0','0'),
            ('1','1','0','1','0','1','1','0','0','1','1','1','1','0'),
            ('1','1','0','1','0','1','1','0','1','0','0','0','0','0'),
            ('1','1','0','1','0','1','1','0','1','0','0','0','1','0'),
            ('1','1','0','1','0','1','1','0','1','0','0','1','0','0'),
            ('1','1','0','1','0','1','1','0','1','0','0','1','1','0'),
            ('1','1','0','1','0','1','1','0','1','0','1','0','0','0'),
            ('1','1','0','1','0','1','1','0','1','0','1','0','1','0'),
            ('1','1','0','1','0','1','1','0','1','0','1','1','0','0'),
            ('1','1','0','1','0','1','1','0','1','0','1','1','1','0'),
            ('1','1','0','1','0','1','1','0','1','1','0','0','0','0'),
            ('1','1','0','1','0','1','1','0','1','1','0','0','1','0'),
            ('1','1','0','1','0','1','1','0','1','1','0','1','0','0'),
            ('1','1','0','1','0','1','1','0','1','1','0','1','1','0'),
            ('1','1','0','1','0','1','1','0','1','1','1','0','0','0'),
            ('1','1','0','1','0','1','1','0','1','1','1','0','1','0'),
            ('1','1','0','1','0','1','1','0','1','1','1','1','0','0'),
            ('1','1','0','1','0','1','1','0','1','1','1','1','1','0'),
            ('1','1','0','1','0','1','1','1','0','0','0','0','0','0'),
            ('1','1','0','1','0','1','1','1','0','0','0','0','1','0'),
            ('1','1','0','1','0','1','1','1','0','0','0','1','0','0'),
            ('1','1','0','1','0','1','1','1','0','0','0','1','1','0'),
            ('1','1','0','1','0','1','1','1','0','0','1','0','0','0'),
            ('1','1','0','1','0','1','1','1','0','0','1','0','1','0'),
            ('1','1','0','1','0','1','1','1','0','0','1','1','0','0'),
            ('1','1','0','1','0','1','1','1','0','0','1','1','1','0'),
            ('1','1','0','1','0','1','1','1','0','1','0','0','0','0'),
            ('1','1','0','1','0','1','1','1','0','1','0','0','1','0'),
            ('1','1','0','1','0','1','1','1','0','1','0','1','0','0'),
            ('1','1','0','1','0','1','1','1','0','1','0','1','1','0'),
            ('1','1','0','1','0','1','1','1','0','1','1','0','0','0'),
            ('1','1','0','1','0','1','1','1','0','1','1','0','1','0'),
            ('1','1','0','1','0','1','1','1','0','1','1','1','0','0'),
            ('1','1','0','1','0','1','1','1','0','1','1','1','1','0'),
            ('1','1','0','1','0','1','1','1','1','0','0','0','0','0'),
            ('1','1','0','1','0','1','1','1','1','0','0','0','1','0'),
            ('1','1','0','1','0','1','1','1','1','0','0','1','0','0'),
            ('1','1','0','1','0','1','1','1','1','0','0','1','1','0'),
            ('1','1','0','1','0','1','1','1','1','0','1','0','0','0'),
            ('1','1','0','1','0','1','1','1','1','0','1','0','1','0'),
            ('1','1','0','1','0','1','1','1','1','0','1','1','0','0'),
            ('1','1','0','1','0','1','1','1','1','0','1','1','1','0'),
            ('1','1','0','1','0','1','1','1','1','1','0','0','0','0'),
            ('1','1','0','1','0','1','1','1','1','1','0','0','1','0'),
            ('1','1','0','1','0','1','1','1','1','1','0','1','0','0'),
            ('1','1','0','1','0','1','1','1','1','1','0','1','1','0'),
            ('1','1','0','1','0','1','1','1','1','1','1','0','0','0'),
            ('1','1','0','1','0','1','1','1','1','1','1','0','1','0'),
            ('1','1','0','1','0','1','1','1','1','1','1','1','0','0'),
            ('1','1','0','1','0','1','1','1','1','1','1','1','1','0'),
            ('1','1','0','1','1','0','0','0','0','0','0','0','0','0'),
            ('1','1','0','1','1','0','0','0','0','0','0','0','1','0'),
            ('1','1','0','1','1','0','0','0','0','0','0','1','0','0'),
            ('1','1','0','1','1','0','0','0','0','0','0','1','1','0'),
            ('1','1','0','1','1','0','0','0','0','0','1','0','0','0'),
            ('1','1','0','1','1','0','0','0','0','0','1','0','1','0'),
            ('1','1','0','1','1','0','0','0','0','0','1','1','0','0'),
            ('1','1','0','1','1','0','0','0','0','0','1','1','1','0'),
            ('1','1','0','1','1','0','0','0','0','1','0','0','0','0'),
            ('1','1','0','1','1','0','0','0','0','1','0','0','1','0'),
            ('1','1','0','1','1','0','0','0','0','1','0','1','0','0'),
            ('1','1','0','1','1','0','0','0','0','1','0','1','1','0'),
            ('1','1','0','1','1','0','0','0','0','1','1','0','0','0'),
            ('1','1','0','1','1','0','0','0','0','1','1','0','1','0'),
            ('1','1','0','1','1','0','0','0','0','1','1','1','0','0'),
            ('1','1','0','1','1','0','0','0','0','1','1','1','1','0'),
            ('1','1','0','1','1','0','0','0','1','0','0','0','0','0'),
            ('1','1','0','1','1','0','0','0','1','0','0','0','1','0'),
            ('1','1','0','1','1','0','0','0','1','0','0','1','0','0'),
            ('1','1','0','1','1','0','0','0','1','0','0','1','1','0'),
            ('1','1','0','1','1','0','0','0','1','0','1','0','0','0'),
            ('1','1','0','1','1','0','0','0','1','0','1','0','1','0'),
            ('1','1','0','1','1','0','0','0','1','0','1','1','0','0'),
            ('1','1','0','1','1','0','0','0','1','0','1','1','1','0'),
            ('1','1','0','1','1','0','0','0','1','1','0','0','0','0'),
            ('1','1','0','1','1','0','0','0','1','1','0','0','1','0'),
            ('1','1','0','1','1','0','0','0','1','1','0','1','0','0'),
            ('1','1','0','1','1','0','0','0','1','1','0','1','1','0'),
            ('1','1','0','1','1','0','0','0','1','1','1','0','0','0'),
            ('1','1','0','1','1','0','0','0','1','1','1','0','1','0'),
            ('1','1','0','1','1','0','0','0','1','1','1','1','0','0'),
            ('1','1','0','1','1','0','0','0','1','1','1','1','1','0'),
            ('1','1','0','1','1','0','0','1','0','0','0','0','0','0'),
            ('1','1','0','1','1','0','0','1','0','0','0','0','1','0'),
            ('1','1','0','1','1','0','0','1','0','0','0','1','0','0'),
            ('1','1','0','1','1','0','0','1','0','0','0','1','1','0'),
            ('1','1','0','1','1','0','0','1','0','0','1','0','0','0'),
            ('1','1','0','1','1','0','0','1','0','0','1','0','1','0'),
            ('1','1','0','1','1','0','0','1','0','0','1','1','0','0'),
            ('1','1','0','1','1','0','0','1','0','0','1','1','1','0'),
            ('1','1','0','1','1','0','0','1','0','1','0','0','0','0'),
            ('1','1','0','1','1','0','0','1','0','1','0','0','1','0'),
            ('1','1','0','1','1','0','0','1','0','1','0','1','0','0'),
            ('1','1','0','1','1','0','0','1','0','1','0','1','1','0'),
            ('1','1','0','1','1','0','0','1','0','1','1','0','0','0'),
            ('1','1','0','1','1','0','0','1','0','1','1','0','1','0'),
            ('1','1','0','1','1','0','0','1','0','1','1','1','0','0'),
            ('1','1','0','1','1','0','0','1','0','1','1','1','1','0'),
            ('1','1','0','1','1','0','0','1','1','0','0','0','0','0'),
            ('1','1','0','1','1','0','0','1','1','0','0','0','1','0'),
            ('1','1','0','1','1','0','0','1','1','0','0','1','0','0'),
            ('1','1','0','1','1','0','0','1','1','0','0','1','1','0'),
            ('1','1','0','1','1','0','0','1','1','0','1','0','0','0'),
            ('1','1','0','1','1','0','0','1','1','0','1','0','1','0'),
            ('1','1','0','1','1','0','0','1','1','0','1','1','0','0'),
            ('1','1','0','1','1','0','0','1','1','0','1','1','1','0'),
            ('1','1','0','1','1','0','0','1','1','1','0','0','0','0'),
            ('1','1','0','1','1','0','0','1','1','1','0','0','1','0'),
            ('1','1','0','1','1','0','0','1','1','1','0','1','0','0'),
            ('1','1','0','1','1','0','0','1','1','1','0','1','1','0'),
            ('1','1','0','1','1','0','0','1','1','1','1','0','0','0'),
            ('1','1','0','1','1','0','0','1','1','1','1','0','1','0'),
            ('1','1','0','1','1','0','0','1','1','1','1','1','0','0'),
            ('1','1','0','1','1','0','0','1','1','1','1','1','1','0'),
            ('1','1','0','1','1','0','1','0','0','0','0','0','0','0'),
            ('1','1','0','1','1','0','1','0','0','0','0','0','1','0'),
            ('1','1','0','1','1','0','1','0','0','0','0','1','0','0'),
            ('1','1','0','1','1','0','1','0','0','0','0','1','1','0'),
            ('1','1','0','1','1','0','1','0','0','0','1','0','0','0'),
            ('1','1','0','1','1','0','1','0','0','0','1','0','1','0'),
            ('1','1','0','1','1','0','1','0','0','0','1','1','0','0'),
            ('1','1','0','1','1','0','1','0','0','0','1','1','1','0'),
            ('1','1','0','1','1','0','1','0','0','1','0','0','0','0'),
            ('1','1','0','1','1','0','1','0','0','1','0','0','1','0'),
            ('1','1','0','1','1','0','1','0','0','1','0','1','0','0'),
            ('1','1','0','1','1','0','1','0','0','1','0','1','1','0'),
            ('1','1','0','1','1','0','1','0','0','1','1','0','0','0'),
            ('1','1','0','1','1','0','1','0','0','1','1','0','1','0'),
            ('1','1','0','1','1','0','1','0','0','1','1','1','0','0'),
            ('1','1','0','1','1','0','1','0','0','1','1','1','1','0'),
            ('1','1','0','1','1','0','1','0','1','0','0','0','0','0'),
            ('1','1','0','1','1','0','1','0','1','0','0','0','1','0'),
            ('1','1','0','1','1','0','1','0','1','0','0','1','0','0'),
            ('1','1','0','1','1','0','1','0','1','0','0','1','1','0'),
            ('1','1','0','1','1','0','1','0','1','0','1','0','0','0'),
            ('1','1','0','1','1','0','1','0','1','0','1','0','1','0'),
            ('1','1','0','1','1','0','1','0','1','0','1','1','0','0'),
            ('1','1','0','1','1','0','1','0','1','0','1','1','1','0'),
            ('1','1','0','1','1','0','1','0','1','1','0','0','0','0'),
            ('1','1','0','1','1','0','1','0','1','1','0','0','1','0'),
            ('1','1','0','1','1','0','1','0','1','1','0','1','0','0'),
            ('1','1','0','1','1','0','1','0','1','1','0','1','1','0'),
            ('1','1','0','1','1','0','1','0','1','1','1','0','0','0'),
            ('1','1','0','1','1','0','1','0','1','1','1','0','1','0'),
            ('1','1','0','1','1','0','1','0','1','1','1','1','0','0'),
            ('1','1','0','1','1','0','1','0','1','1','1','1','1','0'),
            ('1','1','0','1','1','0','1','1','0','0','0','0','0','0'),
            ('1','1','0','1','1','0','1','1','0','0','0','0','1','0'),
            ('1','1','0','1','1','0','1','1','0','0','0','1','0','0'),
            ('1','1','0','1','1','0','1','1','0','0','0','1','1','0'),
            ('1','1','0','1','1','0','1','1','0','0','1','0','0','0'),
            ('1','1','0','1','1','0','1','1','0','0','1','0','1','0'),
            ('1','1','0','1','1','0','1','1','0','0','1','1','0','0'),
            ('1','1','0','1','1','0','1','1','0','0','1','1','1','0'),
            ('1','1','0','1','1','0','1','1','0','1','0','0','0','0'),
            ('1','1','0','1','1','0','1','1','0','1','0','0','1','0'),
            ('1','1','0','1','1','0','1','1','0','1','0','1','0','0'),
            ('1','1','0','1','1','0','1','1','0','1','0','1','1','0'),
            ('1','1','0','1','1','0','1','1','0','1','1','0','0','0'),
            ('1','1','0','1','1','0','1','1','0','1','1','0','1','0'),
            ('1','1','0','1','1','0','1','1','0','1','1','1','0','0'),
            ('1','1','0','1','1','0','1','1','0','1','1','1','1','0'),
            ('1','1','0','1','1','0','1','1','1','0','0','0','0','0'),
            ('1','1','0','1','1','0','1','1','1','0','0','0','1','0'),
            ('1','1','0','1','1','0','1','1','1','0','0','1','0','0'),
            ('1','1','0','1','1','0','1','1','1','0','0','1','1','0'),
            ('1','1','0','1','1','0','1','1','1','0','1','0','0','0'),
            ('1','1','0','1','1','0','1','1','1','0','1','0','1','0'),
            ('1','1','0','1','1','0','1','1','1','0','1','1','0','0'),
            ('1','1','0','1','1','0','1','1','1','0','1','1','1','0'),
            ('1','1','0','1','1','0','1','1','1','1','0','0','0','0'),
            ('1','1','0','1','1','0','1','1','1','1','0','0','1','0'),
            ('1','1','0','1','1','0','1','1','1','1','0','1','0','0'),
            ('1','1','0','1','1','0','1','1','1','1','0','1','1','0'),
            ('1','1','0','1','1','0','1','1','1','1','1','0','0','0'),
            ('1','1','0','1','1','0','1','1','1','1','1','0','1','0'),
            ('1','1','0','1','1','0','1','1','1','1','1','1','0','0'),
            ('1','1','0','1','1','0','1','1','1','1','1','1','1','0'),
            ('1','1','0','1','1','1','0','0','0','0','0','0','0','0'),
            ('1','1','0','1','1','1','0','0','0','0','0','0','1','0'),
            ('1','1','0','1','1','1','0','0','0','0','0','1','0','0'),
            ('1','1','0','1','1','1','0','0','0','0','0','1','1','0'),
            ('1','1','0','1','1','1','0','0','0','0','1','0','0','0'),
            ('1','1','0','1','1','1','0','0','0','0','1','0','1','0'),
            ('1','1','0','1','1','1','0','0','0','0','1','1','0','0'),
            ('1','1','0','1','1','1','0','0','0','0','1','1','1','0'),
            ('1','1','0','1','1','1','0','0','0','1','0','0','0','0'),
            ('1','1','0','1','1','1','0','0','0','1','0','0','1','0'),
            ('1','1','0','1','1','1','0','0','0','1','0','1','0','0'),
            ('1','1','0','1','1','1','0','0','0','1','0','1','1','0'),
            ('1','1','0','1','1','1','0','0','0','1','1','0','0','0'),
            ('1','1','0','1','1','1','0','0','0','1','1','0','1','0'),
            ('1','1','0','1','1','1','0','0','0','1','1','1','0','0'),
            ('1','1','0','1','1','1','0','0','0','1','1','1','1','0'),
            ('1','1','0','1','1','1','0','0','1','0','0','0','0','0'),
            ('1','1','0','1','1','1','0','0','1','0','0','0','1','0'),
            ('1','1','0','1','1','1','0','0','1','0','0','1','0','0'),
            ('1','1','0','1','1','1','0','0','1','0','0','1','1','0'),
            ('1','1','0','1','1','1','0','0','1','0','1','0','0','0'),
            ('1','1','0','1','1','1','0','0','1','0','1','0','1','0'),
            ('1','1','0','1','1','1','0','0','1','0','1','1','0','0'),
            ('1','1','0','1','1','1','0','0','1','0','1','1','1','0'),
            ('1','1','0','1','1','1','0','0','1','1','0','0','0','0'),
            ('1','1','0','1','1','1','0','0','1','1','0','0','1','0'),
            ('1','1','0','1','1','1','0','0','1','1','0','1','0','0'),
            ('1','1','0','1','1','1','0','0','1','1','0','1','1','0'),
            ('1','1','0','1','1','1','0','0','1','1','1','0','0','0'),
            ('1','1','0','1','1','1','0','0','1','1','1','0','1','0'),
            ('1','1','0','1','1','1','0','0','1','1','1','1','0','0'),
            ('1','1','0','1','1','1','0','0','1','1','1','1','1','0'),
            ('1','1','0','1','1','1','0','1','0','0','0','0','0','0'),
            ('1','1','0','1','1','1','0','1','0','0','0','0','1','0'),
            ('1','1','0','1','1','1','0','1','0','0','0','1','0','0'),
            ('1','1','0','1','1','1','0','1','0','0','0','1','1','0'),
            ('1','1','0','1','1','1','0','1','0','0','1','0','0','0'),
            ('1','1','0','1','1','1','0','1','0','0','1','0','1','0'),
            ('1','1','0','1','1','1','0','1','0','0','1','1','0','0'),
            ('1','1','0','1','1','1','0','1','0','0','1','1','1','0'),
            ('1','1','0','1','1','1','0','1','0','1','0','0','0','0'),
            ('1','1','0','1','1','1','0','1','0','1','0','0','1','0'),
            ('1','1','0','1','1','1','0','1','0','1','0','1','0','0'),
            ('1','1','0','1','1','1','0','1','0','1','0','1','1','0'),
            ('1','1','0','1','1','1','0','1','0','1','1','0','0','0'),
            ('1','1','0','1','1','1','0','1','0','1','1','0','1','0'),
            ('1','1','0','1','1','1','0','1','0','1','1','1','0','0'),
            ('1','1','0','1','1','1','0','1','0','1','1','1','1','0'),
            ('1','1','0','1','1','1','0','1','1','0','0','0','0','0'),
            ('1','1','0','1','1','1','0','1','1','0','0','0','1','0'),
            ('1','1','0','1','1','1','0','1','1','0','0','1','0','0'),
            ('1','1','0','1','1','1','0','1','1','0','0','1','1','0'),
            ('1','1','0','1','1','1','0','1','1','0','1','0','0','0'),
            ('1','1','0','1','1','1','0','1','1','0','1','0','1','0'),
            ('1','1','0','1','1','1','0','1','1','0','1','1','0','0'),
            ('1','1','0','1','1','1','0','1','1','0','1','1','1','0'),
            ('1','1','0','1','1','1','0','1','1','1','0','0','0','0'),
            ('1','1','0','1','1','1','0','1','1','1','0','0','1','0'),
            ('1','1','0','1','1','1','0','1','1','1','0','1','0','0'),
            ('1','1','0','1','1','1','0','1','1','1','0','1','1','0'),
            ('1','1','0','1','1','1','0','1','1','1','1','0','0','0'),
            ('1','1','0','1','1','1','0','1','1','1','1','0','1','0'),
            ('1','1','0','1','1','1','0','1','1','1','1','1','0','0'),
            ('1','1','0','1','1','1','0','1','1','1','1','1','1','0'),
            ('1','1','0','1','1','1','1','0','0','0','0','0','0','0'),
            ('1','1','0','1','1','1','1','0','0','0','0','0','1','0'),
            ('1','1','0','1','1','1','1','0','0','0','0','1','0','0'),
            ('1','1','0','1','1','1','1','0','0','0','0','1','1','0'),
            ('1','1','0','1','1','1','1','0','0','0','1','0','0','0'),
            ('1','1','0','1','1','1','1','0','0','0','1','0','1','0'),
            ('1','1','0','1','1','1','1','0','0','0','1','1','0','0'),
            ('1','1','0','1','1','1','1','0','0','0','1','1','1','0'),
            ('1','1','0','1','1','1','1','0','0','1','0','0','0','0'),
            ('1','1','0','1','1','1','1','0','0','1','0','0','1','0'),
            ('1','1','0','1','1','1','1','0','0','1','0','1','0','0'),
            ('1','1','0','1','1','1','1','0','0','1','0','1','1','0'),
            ('1','1','0','1','1','1','1','0','0','1','1','0','0','0'),
            ('1','1','0','1','1','1','1','0','0','1','1','0','1','0'),
            ('1','1','0','1','1','1','1','0','0','1','1','1','0','0'),
            ('1','1','0','1','1','1','1','0','0','1','1','1','1','0'),
            ('1','1','0','1','1','1','1','0','1','0','0','0','0','0'),
            ('1','1','0','1','1','1','1','0','1','0','0','0','1','0'),
            ('1','1','0','1','1','1','1','0','1','0','0','1','0','0'),
            ('1','1','0','1','1','1','1','0','1','0','0','1','1','0'),
            ('1','1','0','1','1','1','1','0','1','0','1','0','0','0'),
            ('1','1','0','1','1','1','1','0','1','0','1','0','1','0'),
            ('1','1','0','1','1','1','1','0','1','0','1','1','0','0'),
            ('1','1','0','1','1','1','1','0','1','0','1','1','1','0'),
            ('1','1','0','1','1','1','1','0','1','1','0','0','0','0'),
            ('1','1','0','1','1','1','1','0','1','1','0','0','1','0'),
            ('1','1','0','1','1','1','1','0','1','1','0','1','0','0'),
            ('1','1','0','1','1','1','1','0','1','1','0','1','1','0'),
            ('1','1','0','1','1','1','1','0','1','1','1','0','0','0'),
            ('1','1','0','1','1','1','1','0','1','1','1','0','1','0'),
            ('1','1','0','1','1','1','1','0','1','1','1','1','0','0'),
            ('1','1','0','1','1','1','1','0','1','1','1','1','1','0'),
            ('1','1','0','1','1','1','1','1','0','0','0','0','0','0'),
            ('1','1','0','1','1','1','1','1','0','0','0','0','1','0'),
            ('1','1','0','1','1','1','1','1','0','0','0','1','0','0'),
            ('1','1','0','1','1','1','1','1','0','0','0','1','1','0'),
            ('1','1','0','1','1','1','1','1','0','0','1','0','0','0'),
            ('1','1','0','1','1','1','1','1','0','0','1','0','1','0'),
            ('1','1','0','1','1','1','1','1','0','0','1','1','0','0'),
            ('1','1','0','1','1','1','1','1','0','0','1','1','1','0'),
            ('1','1','0','1','1','1','1','1','0','1','0','0','0','0'),
            ('1','1','0','1','1','1','1','1','0','1','0','0','1','0'),
            ('1','1','0','1','1','1','1','1','0','1','0','1','0','0'),
            ('1','1','0','1','1','1','1','1','0','1','0','1','1','0'),
            ('1','1','0','1','1','1','1','1','0','1','1','0','0','0'),
            ('1','1','0','1','1','1','1','1','0','1','1','0','1','0'),
            ('1','1','0','1','1','1','1','1','0','1','1','1','0','0'),
            ('1','1','0','1','1','1','1','1','0','1','1','1','1','0'),
            ('1','1','0','1','1','1','1','1','1','0','0','0','0','0'),
            ('1','1','0','1','1','1','1','1','1','0','0','0','1','0'),
            ('1','1','0','1','1','1','1','1','1','0','0','1','0','0'),
            ('1','1','0','1','1','1','1','1','1','0','0','1','1','0'),
            ('1','1','0','1','1','1','1','1','1','0','1','0','0','0'),
            ('1','1','0','1','1','1','1','1','1','0','1','0','1','0'),
            ('1','1','0','1','1','1','1','1','1','0','1','1','0','0'),
            ('1','1','0','1','1','1','1','1','1','0','1','1','1','0'),
            ('1','1','0','1','1','1','1','1','1','1','0','0','0','0'),
            ('1','1','0','1','1','1','1','1','1','1','0','0','1','0'),
            ('1','1','0','1','1','1','1','1','1','1','0','1','0','0'),
            ('1','1','0','1','1','1','1','1','1','1','0','1','1','0'),
            ('1','1','0','1','1','1','1','1','1','1','1','0','0','0'),
            ('1','1','0','1','1','1','1','1','1','1','1','0','1','0'),
            ('1','1','0','1','1','1','1','1','1','1','1','1','0','0'),
            ('1','1','0','1','1','1','1','1','1','1','1','1','1','0'),
            ('1','1','1','0','0','0','0','0','0','0','0','0','0','0'),
            ('1','1','1','0','0','0','0','0','0','0','0','0','1','0'),
            ('1','1','1','0','0','0','0','0','0','0','0','1','0','0'),
            ('1','1','1','0','0','0','0','0','0','0','0','1','1','0'),
            ('1','1','1','0','0','0','0','0','0','0','1','0','0','0'),
            ('1','1','1','0','0','0','0','0','0','0','1','0','1','0'),
            ('1','1','1','0','0','0','0','0','0','0','1','1','0','0'),
            ('1','1','1','0','0','0','0','0','0','0','1','1','1','0'),
            ('1','1','1','0','0','0','0','0','0','1','0','0','0','0'),
            ('1','1','1','0','0','0','0','0','0','1','0','0','1','0'),
            ('1','1','1','0','0','0','0','0','0','1','0','1','0','0'),
            ('1','1','1','0','0','0','0','0','0','1','0','1','1','0'),
            ('1','1','1','0','0','0','0','0','0','1','1','0','0','0'),
            ('1','1','1','0','0','0','0','0','0','1','1','0','1','0'),
            ('1','1','1','0','0','0','0','0','0','1','1','1','0','0'),
            ('1','1','1','0','0','0','0','0','0','1','1','1','1','0'),
            ('1','1','1','0','0','0','0','0','1','0','0','0','0','0'),
            ('1','1','1','0','0','0','0','0','1','0','0','0','1','0'),
            ('1','1','1','0','0','0','0','0','1','0','0','1','0','0'),
            ('1','1','1','0','0','0','0','0','1','0','0','1','1','0'),
            ('1','1','1','0','0','0','0','0','1','0','1','0','0','0'),
            ('1','1','1','0','0','0','0','0','1','0','1','0','1','0'),
            ('1','1','1','0','0','0','0','0','1','0','1','1','0','0'),
            ('1','1','1','0','0','0','0','0','1','0','1','1','1','0'),
            ('1','1','1','0','0','0','0','0','1','1','0','0','0','0'),
            ('1','1','1','0','0','0','0','0','1','1','0','0','1','0'),
            ('1','1','1','0','0','0','0','0','1','1','0','1','0','0'),
            ('1','1','1','0','0','0','0','0','1','1','0','1','1','0'),
            ('1','1','1','0','0','0','0','0','1','1','1','0','0','0'),
            ('1','1','1','0','0','0','0','0','1','1','1','0','1','0'),
            ('1','1','1','0','0','0','0','0','1','1','1','1','0','0'),
            ('1','1','1','0','0','0','0','0','1','1','1','1','1','0'),
            ('1','1','1','0','0','0','0','1','0','0','0','0','0','0'),
            ('1','1','1','0','0','0','0','1','0','0','0','0','1','0'),
            ('1','1','1','0','0','0','0','1','0','0','0','1','0','0'),
            ('1','1','1','0','0','0','0','1','0','0','0','1','1','0'),
            ('1','1','1','0','0','0','0','1','0','0','1','0','0','0'),
            ('1','1','1','0','0','0','0','1','0','0','1','0','1','0'),
            ('1','1','1','0','0','0','0','1','0','0','1','1','0','0'),
            ('1','1','1','0','0','0','0','1','0','0','1','1','1','0'),
            ('1','1','1','0','0','0','0','1','0','1','0','0','0','0'),
            ('1','1','1','0','0','0','0','1','0','1','0','0','1','0'),
            ('1','1','1','0','0','0','0','1','0','1','0','1','0','0'),
            ('1','1','1','0','0','0','0','1','0','1','0','1','1','0'),
            ('1','1','1','0','0','0','0','1','0','1','1','0','0','0'),
            ('1','1','1','0','0','0','0','1','0','1','1','0','1','0'),
            ('1','1','1','0','0','0','0','1','0','1','1','1','0','0'),
            ('1','1','1','0','0','0','0','1','0','1','1','1','1','0'),
            ('1','1','1','0','0','0','0','1','1','0','0','0','0','0'),
            ('1','1','1','0','0','0','0','1','1','0','0','0','1','0'),
            ('1','1','1','0','0','0','0','1','1','0','0','1','0','0'),
            ('1','1','1','0','0','0','0','1','1','0','0','1','1','0'),
            ('1','1','1','0','0','0','0','1','1','0','1','0','0','0'),
            ('1','1','1','0','0','0','0','1','1','0','1','0','1','0'),
            ('1','1','1','0','0','0','0','1','1','0','1','1','0','0'),
            ('1','1','1','0','0','0','0','1','1','0','1','1','1','0'),
            ('1','1','1','0','0','0','0','1','1','1','0','0','0','0'),
            ('1','1','1','0','0','0','0','1','1','1','0','0','1','0'),
            ('1','1','1','0','0','0','0','1','1','1','0','1','0','0'),
            ('1','1','1','0','0','0','0','1','1','1','0','1','1','0'),
            ('1','1','1','0','0','0','0','1','1','1','1','0','0','0'),
            ('1','1','1','0','0','0','0','1','1','1','1','0','1','0'),
            ('1','1','1','0','0','0','0','1','1','1','1','1','0','0'),
            ('1','1','1','0','0','0','0','1','1','1','1','1','1','0'),
            ('1','1','1','0','0','0','1','0','0','0','0','0','0','0'),
            ('1','1','1','0','0','0','1','0','0','0','0','0','1','0'),
            ('1','1','1','0','0','0','1','0','0','0','0','1','0','0'),
            ('1','1','1','0','0','0','1','0','0','0','0','1','1','0'),
            ('1','1','1','0','0','0','1','0','0','0','1','0','0','0'),
            ('1','1','1','0','0','0','1','0','0','0','1','0','1','0'),
            ('1','1','1','0','0','0','1','0','0','0','1','1','0','0'),
            ('1','1','1','0','0','0','1','0','0','0','1','1','1','0'),
            ('1','1','1','0','0','0','1','0','0','1','0','0','0','0'),
            ('1','1','1','0','0','0','1','0','0','1','0','0','1','0'),
            ('1','1','1','0','0','0','1','0','0','1','0','1','0','0'),
            ('1','1','1','0','0','0','1','0','0','1','0','1','1','0'),
            ('1','1','1','0','0','0','1','0','0','1','1','0','0','0'),
            ('1','1','1','0','0','0','1','0','0','1','1','0','1','0'),
            ('1','1','1','0','0','0','1','0','0','1','1','1','0','0'),
            ('1','1','1','0','0','0','1','0','0','1','1','1','1','0'),
            ('1','1','1','0','0','0','1','0','1','0','0','0','0','0'),
            ('1','1','1','0','0','0','1','0','1','0','0','0','1','0'),
            ('1','1','1','0','0','0','1','0','1','0','0','1','0','0'),
            ('1','1','1','0','0','0','1','0','1','0','0','1','1','0'),
            ('1','1','1','0','0','0','1','0','1','0','1','0','0','0'),
            ('1','1','1','0','0','0','1','0','1','0','1','0','1','0'),
            ('1','1','1','0','0','0','1','0','1','0','1','1','0','0'),
            ('1','1','1','0','0','0','1','0','1','0','1','1','1','0'),
            ('1','1','1','0','0','0','1','0','1','1','0','0','0','0'),
            ('1','1','1','0','0','0','1','0','1','1','0','0','1','0'),
            ('1','1','1','0','0','0','1','0','1','1','0','1','0','0'),
            ('1','1','1','0','0','0','1','0','1','1','0','1','1','0'),
            ('1','1','1','0','0','0','1','0','1','1','1','0','0','0'),
            ('1','1','1','0','0','0','1','0','1','1','1','0','1','0'),
            ('1','1','1','0','0','0','1','0','1','1','1','1','0','0'),
            ('1','1','1','0','0','0','1','0','1','1','1','1','1','0'),
            ('1','1','1','0','0','0','1','1','0','0','0','0','0','0'),
            ('1','1','1','0','0','0','1','1','0','0','0','0','1','0'),
            ('1','1','1','0','0','0','1','1','0','0','0','1','0','0'),
            ('1','1','1','0','0','0','1','1','0','0','0','1','1','0'),
            ('1','1','1','0','0','0','1','1','0','0','1','0','0','0'),
            ('1','1','1','0','0','0','1','1','0','0','1','0','1','0'),
            ('1','1','1','0','0','0','1','1','0','0','1','1','0','0'),
            ('1','1','1','0','0','0','1','1','0','0','1','1','1','0'),
            ('1','1','1','0','0','0','1','1','0','1','0','0','0','0'),
            ('1','1','1','0','0','0','1','1','0','1','0','0','1','0'),
            ('1','1','1','0','0','0','1','1','0','1','0','1','0','0'),
            ('1','1','1','0','0','0','1','1','0','1','0','1','1','0'),
            ('1','1','1','0','0','0','1','1','0','1','1','0','0','0'),
            ('1','1','1','0','0','0','1','1','0','1','1','0','1','0'),
            ('1','1','1','0','0','0','1','1','0','1','1','1','0','0'),
            ('1','1','1','0','0','0','1','1','0','1','1','1','1','0'),
            ('1','1','1','0','0','0','1','1','1','0','0','0','0','0'),
            ('1','1','1','0','0','0','1','1','1','0','0','0','1','0'),
            ('1','1','1','0','0','0','1','1','1','0','0','1','0','0'),
            ('1','1','1','0','0','0','1','1','1','0','0','1','1','0'),
            ('1','1','1','0','0','0','1','1','1','0','1','0','0','0'),
            ('1','1','1','0','0','0','1','1','1','0','1','0','1','0'),
            ('1','1','1','0','0','0','1','1','1','0','1','1','0','0'),
            ('1','1','1','0','0','0','1','1','1','0','1','1','1','0'),
            ('1','1','1','0','0','0','1','1','1','1','0','0','0','0'),
            ('1','1','1','0','0','0','1','1','1','1','0','0','1','0'),
            ('1','1','1','0','0','0','1','1','1','1','0','1','0','0'),
            ('1','1','1','0','0','0','1','1','1','1','0','1','1','0'),
            ('1','1','1','0','0','0','1','1','1','1','1','0','0','0'),
            ('1','1','1','0','0','0','1','1','1','1','1','0','1','0'),
            ('1','1','1','0','0','0','1','1','1','1','1','1','0','0'),
            ('1','1','1','0','0','0','1','1','1','1','1','1','1','0'),
            ('1','1','1','0','0','1','0','0','0','0','0','0','0','0'),
            ('1','1','1','0','0','1','0','0','0','0','0','0','1','0'),
            ('1','1','1','0','0','1','0','0','0','0','0','1','0','0'),
            ('1','1','1','0','0','1','0','0','0','0','0','1','1','0'),
            ('1','1','1','0','0','1','0','0','0','0','1','0','0','0'),
            ('1','1','1','0','0','1','0','0','0','0','1','0','1','0'),
            ('1','1','1','0','0','1','0','0','0','0','1','1','0','0'),
            ('1','1','1','0','0','1','0','0','0','0','1','1','1','0'),
            ('1','1','1','0','0','1','0','0','0','1','0','0','0','0'),
            ('1','1','1','0','0','1','0','0','0','1','0','0','1','0'),
            ('1','1','1','0','0','1','0','0','0','1','0','1','0','0'),
            ('1','1','1','0','0','1','0','0','0','1','0','1','1','0'),
            ('1','1','1','0','0','1','0','0','0','1','1','0','0','0'),
            ('1','1','1','0','0','1','0','0','0','1','1','0','1','0'),
            ('1','1','1','0','0','1','0','0','0','1','1','1','0','0'),
            ('1','1','1','0','0','1','0','0','0','1','1','1','1','0'),
            ('1','1','1','0','0','1','0','0','1','0','0','0','0','0'),
            ('1','1','1','0','0','1','0','0','1','0','0','0','1','0'),
            ('1','1','1','0','0','1','0','0','1','0','0','1','0','0'),
            ('1','1','1','0','0','1','0','0','1','0','0','1','1','0'),
            ('1','1','1','0','0','1','0','0','1','0','1','0','0','0'),
            ('1','1','1','0','0','1','0','0','1','0','1','0','1','0'),
            ('1','1','1','0','0','1','0','0','1','0','1','1','0','0'),
            ('1','1','1','0','0','1','0','0','1','0','1','1','1','0'),
            ('1','1','1','0','0','1','0','0','1','1','0','0','0','0'),
            ('1','1','1','0','0','1','0','0','1','1','0','0','1','0'),
            ('1','1','1','0','0','1','0','0','1','1','0','1','0','0'),
            ('1','1','1','0','0','1','0','0','1','1','0','1','1','0'),
            ('1','1','1','0','0','1','0','0','1','1','1','0','0','0'),
            ('1','1','1','0','0','1','0','0','1','1','1','0','1','0'),
            ('1','1','1','0','0','1','0','0','1','1','1','1','0','0'),
            ('1','1','1','0','0','1','0','0','1','1','1','1','1','0'),
            ('1','1','1','0','0','1','0','1','0','0','0','0','0','0'),
            ('1','1','1','0','0','1','0','1','0','0','0','0','1','0'),
            ('1','1','1','0','0','1','0','1','0','0','0','1','0','0'),
            ('1','1','1','0','0','1','0','1','0','0','0','1','1','0'),
            ('1','1','1','0','0','1','0','1','0','0','1','0','0','0'),
            ('1','1','1','0','0','1','0','1','0','0','1','0','1','0'),
            ('1','1','1','0','0','1','0','1','0','0','1','1','0','0'),
            ('1','1','1','0','0','1','0','1','0','0','1','1','1','0'),
            ('1','1','1','0','0','1','0','1','0','1','0','0','0','0'),
            ('1','1','1','0','0','1','0','1','0','1','0','0','1','0'),
            ('1','1','1','0','0','1','0','1','0','1','0','1','0','0'),
            ('1','1','1','0','0','1','0','1','0','1','0','1','1','0'),
            ('1','1','1','0','0','1','0','1','0','1','1','0','0','0'),
            ('1','1','1','0','0','1','0','1','0','1','1','0','1','0'),
            ('1','1','1','0','0','1','0','1','0','1','1','1','0','0'),
            ('1','1','1','0','0','1','0','1','0','1','1','1','1','0'),
            ('1','1','1','0','0','1','0','1','1','0','0','0','0','0'),
            ('1','1','1','0','0','1','0','1','1','0','0','0','1','0'),
            ('1','1','1','0','0','1','0','1','1','0','0','1','0','0'),
            ('1','1','1','0','0','1','0','1','1','0','0','1','1','0'),
            ('1','1','1','0','0','1','0','1','1','0','1','0','0','0'),
            ('1','1','1','0','0','1','0','1','1','0','1','0','1','0'),
            ('1','1','1','0','0','1','0','1','1','0','1','1','0','0'),
            ('1','1','1','0','0','1','0','1','1','0','1','1','1','0'),
            ('1','1','1','0','0','1','0','1','1','1','0','0','0','0'),
            ('1','1','1','0','0','1','0','1','1','1','0','0','1','0'),
            ('1','1','1','0','0','1','0','1','1','1','0','1','0','0'),
            ('1','1','1','0','0','1','0','1','1','1','0','1','1','0'),
            ('1','1','1','0','0','1','0','1','1','1','1','0','0','0'),
            ('1','1','1','0','0','1','0','1','1','1','1','0','1','0'),
            ('1','1','1','0','0','1','0','1','1','1','1','1','0','0'),
            ('1','1','1','0','0','1','0','1','1','1','1','1','1','0'),
            ('1','1','1','0','0','1','1','0','0','0','0','0','0','0'),
            ('1','1','1','0','0','1','1','0','0','0','0','0','1','0'),
            ('1','1','1','0','0','1','1','0','0','0','0','1','0','0'),
            ('1','1','1','0','0','1','1','0','0','0','0','1','1','0'),
            ('1','1','1','0','0','1','1','0','0','0','1','0','0','0'),
            ('1','1','1','0','0','1','1','0','0','0','1','0','1','0'),
            ('1','1','1','0','0','1','1','0','0','0','1','1','0','0'),
            ('1','1','1','0','0','1','1','0','0','0','1','1','1','0'),
            ('1','1','1','0','0','1','1','0','0','1','0','0','0','0'),
            ('1','1','1','0','0','1','1','0','0','1','0','0','1','0'),
            ('1','1','1','0','0','1','1','0','0','1','0','1','0','0'),
            ('1','1','1','0','0','1','1','0','0','1','0','1','1','0'),
            ('1','1','1','0','0','1','1','0','0','1','1','0','0','0'),
            ('1','1','1','0','0','1','1','0','0','1','1','0','1','0'),
            ('1','1','1','0','0','1','1','0','0','1','1','1','0','0'),
            ('1','1','1','0','0','1','1','0','0','1','1','1','1','0'),
            ('1','1','1','0','0','1','1','0','1','0','0','0','0','0'),
            ('1','1','1','0','0','1','1','0','1','0','0','0','1','0'),
            ('1','1','1','0','0','1','1','0','1','0','0','1','0','0'),
            ('1','1','1','0','0','1','1','0','1','0','0','1','1','0'),
            ('1','1','1','0','0','1','1','0','1','0','1','0','0','0'),
            ('1','1','1','0','0','1','1','0','1','0','1','0','1','0'),
            ('1','1','1','0','0','1','1','0','1','0','1','1','0','0'),
            ('1','1','1','0','0','1','1','0','1','0','1','1','1','0'),
            ('1','1','1','0','0','1','1','0','1','1','0','0','0','0'),
            ('1','1','1','0','0','1','1','0','1','1','0','0','1','0'),
            ('1','1','1','0','0','1','1','0','1','1','0','1','0','0'),
            ('1','1','1','0','0','1','1','0','1','1','0','1','1','0'),
            ('1','1','1','0','0','1','1','0','1','1','1','0','0','0'),
            ('1','1','1','0','0','1','1','0','1','1','1','0','1','0'),
            ('1','1','1','0','0','1','1','0','1','1','1','1','0','0'),
            ('1','1','1','0','0','1','1','0','1','1','1','1','1','0'),
            ('1','1','1','0','0','1','1','1','0','0','0','0','0','0'),
            ('1','1','1','0','0','1','1','1','0','0','0','0','1','0'),
            ('1','1','1','0','0','1','1','1','0','0','0','1','0','0'),
            ('1','1','1','0','0','1','1','1','0','0','0','1','1','0'),
            ('1','1','1','0','0','1','1','1','0','0','1','0','0','0'),
            ('1','1','1','0','0','1','1','1','0','0','1','0','1','0'),
            ('1','1','1','0','0','1','1','1','0','0','1','1','0','0'),
            ('1','1','1','0','0','1','1','1','0','0','1','1','1','0'),
            ('1','1','1','0','0','1','1','1','0','1','0','0','0','0'),
            ('1','1','1','0','0','1','1','1','0','1','0','0','1','0'),
            ('1','1','1','0','0','1','1','1','0','1','0','1','0','0'),
            ('1','1','1','0','0','1','1','1','0','1','0','1','1','0'),
            ('1','1','1','0','0','1','1','1','0','1','1','0','0','0'),
            ('1','1','1','0','0','1','1','1','0','1','1','0','1','0'),
            ('1','1','1','0','0','1','1','1','0','1','1','1','0','0'),
            ('1','1','1','0','0','1','1','1','0','1','1','1','1','0'),
            ('1','1','1','0','0','1','1','1','1','0','0','0','0','0'),
            ('1','1','1','0','0','1','1','1','1','0','0','0','1','0'),
            ('1','1','1','0','0','1','1','1','1','0','0','1','0','0'),
            ('1','1','1','0','0','1','1','1','1','0','0','1','1','0'),
            ('1','1','1','0','0','1','1','1','1','0','1','0','0','0'),
            ('1','1','1','0','0','1','1','1','1','0','1','0','1','0'),
            ('1','1','1','0','0','1','1','1','1','0','1','1','0','0'),
            ('1','1','1','0','0','1','1','1','1','0','1','1','1','0'),
            ('1','1','1','0','0','1','1','1','1','1','0','0','0','0'),
            ('1','1','1','0','0','1','1','1','1','1','0','0','1','0'),
            ('1','1','1','0','0','1','1','1','1','1','0','1','0','0'),
            ('1','1','1','0','0','1','1','1','1','1','0','1','1','0'),
            ('1','1','1','0','0','1','1','1','1','1','1','0','0','0'),
            ('1','1','1','0','0','1','1','1','1','1','1','0','1','0'),
            ('1','1','1','0','0','1','1','1','1','1','1','1','0','0'),
            ('1','1','1','0','0','1','1','1','1','1','1','1','1','0'),
            ('1','1','1','0','1','0','0','0','0','0','0','0','0','0'),
            ('1','1','1','0','1','0','0','0','0','0','0','0','1','0'),
            ('1','1','1','0','1','0','0','0','0','0','0','1','0','0'),
            ('1','1','1','0','1','0','0','0','0','0','0','1','1','0'),
            ('1','1','1','0','1','0','0','0','0','0','1','0','0','0'),
            ('1','1','1','0','1','0','0','0','0','0','1','0','1','0'),
            ('1','1','1','0','1','0','0','0','0','0','1','1','0','0'),
            ('1','1','1','0','1','0','0','0','0','0','1','1','1','0'),
            ('1','1','1','0','1','0','0','0','0','1','0','0','0','0'),
            ('1','1','1','0','1','0','0','0','0','1','0','0','1','0'),
            ('1','1','1','0','1','0','0','0','0','1','0','1','0','0'),
            ('1','1','1','0','1','0','0','0','0','1','0','1','1','0'),
            ('1','1','1','0','1','0','0','0','0','1','1','0','0','0'),
            ('1','1','1','0','1','0','0','0','0','1','1','0','1','0'),
            ('1','1','1','0','1','0','0','0','0','1','1','1','0','0'),
            ('1','1','1','0','1','0','0','0','0','1','1','1','1','0'),
            ('1','1','1','0','1','0','0','0','1','0','0','0','0','0'),
            ('1','1','1','0','1','0','0','0','1','0','0','0','1','0'),
            ('1','1','1','0','1','0','0','0','1','0','0','1','0','0'),
            ('1','1','1','0','1','0','0','0','1','0','0','1','1','0'),
            ('1','1','1','0','1','0','0','0','1','0','1','0','0','0'),
            ('1','1','1','0','1','0','0','0','1','0','1','0','1','0'),
            ('1','1','1','0','1','0','0','0','1','0','1','1','0','0'),
            ('1','1','1','0','1','0','0','0','1','0','1','1','1','0'),
            ('1','1','1','0','1','0','0','0','1','1','0','0','0','0'),
            ('1','1','1','0','1','0','0','0','1','1','0','0','1','0'),
            ('1','1','1','0','1','0','0','0','1','1','0','1','0','0'),
            ('1','1','1','0','1','0','0','0','1','1','0','1','1','0'),
            ('1','1','1','0','1','0','0','0','1','1','1','0','0','0'),
            ('1','1','1','0','1','0','0','0','1','1','1','0','1','0'),
            ('1','1','1','0','1','0','0','0','1','1','1','1','0','0'),
            ('1','1','1','0','1','0','0','0','1','1','1','1','1','0'),
            ('1','1','1','0','1','0','0','1','0','0','0','0','0','0'),
            ('1','1','1','0','1','0','0','1','0','0','0','0','1','0'),
            ('1','1','1','0','1','0','0','1','0','0','0','1','0','0'),
            ('1','1','1','0','1','0','0','1','0','0','0','1','1','0'),
            ('1','1','1','0','1','0','0','1','0','0','1','0','0','0'),
            ('1','1','1','0','1','0','0','1','0','0','1','0','1','0'),
            ('1','1','1','0','1','0','0','1','0','0','1','1','0','0'),
            ('1','1','1','0','1','0','0','1','0','0','1','1','1','0'),
            ('1','1','1','0','1','0','0','1','0','1','0','0','0','0'),
            ('1','1','1','0','1','0','0','1','0','1','0','0','1','0'),
            ('1','1','1','0','1','0','0','1','0','1','0','1','0','0'),
            ('1','1','1','0','1','0','0','1','0','1','0','1','1','0'),
            ('1','1','1','0','1','0','0','1','0','1','1','0','0','0'),
            ('1','1','1','0','1','0','0','1','0','1','1','0','1','0'),
            ('1','1','1','0','1','0','0','1','0','1','1','1','0','0'),
            ('1','1','1','0','1','0','0','1','0','1','1','1','1','0'),
            ('1','1','1','0','1','0','0','1','1','0','0','0','0','0'),
            ('1','1','1','0','1','0','0','1','1','0','0','0','1','0'),
            ('1','1','1','0','1','0','0','1','1','0','0','1','0','0'),
            ('1','1','1','0','1','0','0','1','1','0','0','1','1','0'),
            ('1','1','1','0','1','0','0','1','1','0','1','0','0','0'),
            ('1','1','1','0','1','0','0','1','1','0','1','0','1','0'),
            ('1','1','1','0','1','0','0','1','1','0','1','1','0','0'),
            ('1','1','1','0','1','0','0','1','1','0','1','1','1','0'),
            ('1','1','1','0','1','0','0','1','1','1','0','0','0','0'),
            ('1','1','1','0','1','0','0','1','1','1','0','0','1','0'),
            ('1','1','1','0','1','0','0','1','1','1','0','1','0','0'),
            ('1','1','1','0','1','0','0','1','1','1','0','1','1','0'),
            ('1','1','1','0','1','0','0','1','1','1','1','0','0','0'),
            ('1','1','1','0','1','0','0','1','1','1','1','0','1','0'),
            ('1','1','1','0','1','0','0','1','1','1','1','1','0','0'),
            ('1','1','1','0','1','0','0','1','1','1','1','1','1','0'),
            ('1','1','1','0','1','0','1','0','0','0','0','0','0','0'),
            ('1','1','1','0','1','0','1','0','0','0','0','0','1','0'),
            ('1','1','1','0','1','0','1','0','0','0','0','1','0','0'),
            ('1','1','1','0','1','0','1','0','0','0','0','1','1','0'),
            ('1','1','1','0','1','0','1','0','0','0','1','0','0','0'),
            ('1','1','1','0','1','0','1','0','0','0','1','0','1','0'),
            ('1','1','1','0','1','0','1','0','0','0','1','1','0','0'),
            ('1','1','1','0','1','0','1','0','0','0','1','1','1','0'),
            ('1','1','1','0','1','0','1','0','0','1','0','0','0','0'),
            ('1','1','1','0','1','0','1','0','0','1','0','0','1','0'),
            ('1','1','1','0','1','0','1','0','0','1','0','1','0','0'),
            ('1','1','1','0','1','0','1','0','0','1','0','1','1','0'),
            ('1','1','1','0','1','0','1','0','0','1','1','0','0','0'),
            ('1','1','1','0','1','0','1','0','0','1','1','0','1','0'),
            ('1','1','1','0','1','0','1','0','0','1','1','1','0','0'),
            ('1','1','1','0','1','0','1','0','0','1','1','1','1','0'),
            ('1','1','1','0','1','0','1','0','1','0','0','0','0','0'),
            ('1','1','1','0','1','0','1','0','1','0','0','0','1','0'),
            ('1','1','1','0','1','0','1','0','1','0','0','1','0','0'),
            ('1','1','1','0','1','0','1','0','1','0','0','1','1','0'),
            ('1','1','1','0','1','0','1','0','1','0','1','0','0','0'),
            ('1','1','1','0','1','0','1','0','1','0','1','0','1','0'),
            ('1','1','1','0','1','0','1','0','1','0','1','1','0','0'),
            ('1','1','1','0','1','0','1','0','1','0','1','1','1','0'),
            ('1','1','1','0','1','0','1','0','1','1','0','0','0','0'),
            ('1','1','1','0','1','0','1','0','1','1','0','0','1','0'),
            ('1','1','1','0','1','0','1','0','1','1','0','1','0','0'),
            ('1','1','1','0','1','0','1','0','1','1','0','1','1','0'),
            ('1','1','1','0','1','0','1','0','1','1','1','0','0','0'),
            ('1','1','1','0','1','0','1','0','1','1','1','0','1','0'),
            ('1','1','1','0','1','0','1','0','1','1','1','1','0','0'),
            ('1','1','1','0','1','0','1','0','1','1','1','1','1','0'),
            ('1','1','1','0','1','0','1','1','0','0','0','0','0','0'),
            ('1','1','1','0','1','0','1','1','0','0','0','0','1','0'),
            ('1','1','1','0','1','0','1','1','0','0','0','1','0','0'),
            ('1','1','1','0','1','0','1','1','0','0','0','1','1','0'),
            ('1','1','1','0','1','0','1','1','0','0','1','0','0','0'),
            ('1','1','1','0','1','0','1','1','0','0','1','0','1','0'),
            ('1','1','1','0','1','0','1','1','0','0','1','1','0','0'),
            ('1','1','1','0','1','0','1','1','0','0','1','1','1','0'),
            ('1','1','1','0','1','0','1','1','0','1','0','0','0','0'),
            ('1','1','1','0','1','0','1','1','0','1','0','0','1','0'),
            ('1','1','1','0','1','0','1','1','0','1','0','1','0','0'),
            ('1','1','1','0','1','0','1','1','0','1','0','1','1','0'),
            ('1','1','1','0','1','0','1','1','0','1','1','0','0','0'),
            ('1','1','1','0','1','0','1','1','0','1','1','0','1','0'),
            ('1','1','1','0','1','0','1','1','0','1','1','1','0','0'),
            ('1','1','1','0','1','0','1','1','0','1','1','1','1','0'),
            ('1','1','1','0','1','0','1','1','1','0','0','0','0','0'),
            ('1','1','1','0','1','0','1','1','1','0','0','0','1','0'),
            ('1','1','1','0','1','0','1','1','1','0','0','1','0','0'),
            ('1','1','1','0','1','0','1','1','1','0','0','1','1','0'),
            ('1','1','1','0','1','0','1','1','1','0','1','0','0','0'),
            ('1','1','1','0','1','0','1','1','1','0','1','0','1','0'),
            ('1','1','1','0','1','0','1','1','1','0','1','1','0','0'),
            ('1','1','1','0','1','0','1','1','1','0','1','1','1','0'),
            ('1','1','1','0','1','0','1','1','1','1','0','0','0','0'),
            ('1','1','1','0','1','0','1','1','1','1','0','0','1','0'),
            ('1','1','1','0','1','0','1','1','1','1','0','1','0','0'),
            ('1','1','1','0','1','0','1','1','1','1','0','1','1','0'),
            ('1','1','1','0','1','0','1','1','1','1','1','0','0','0'),
            ('1','1','1','0','1','0','1','1','1','1','1','0','1','0'),
            ('1','1','1','0','1','0','1','1','1','1','1','1','0','0'),
            ('1','1','1','0','1','0','1','1','1','1','1','1','1','0'),
            ('1','1','1','0','1','1','0','0','0','0','0','0','0','0'),
            ('1','1','1','0','1','1','0','0','0','0','0','0','1','0'),
            ('1','1','1','0','1','1','0','0','0','0','0','1','0','0'),
            ('1','1','1','0','1','1','0','0','0','0','0','1','1','0'),
            ('1','1','1','0','1','1','0','0','0','0','1','0','0','0'),
            ('1','1','1','0','1','1','0','0','0','0','1','0','1','0'),
            ('1','1','1','0','1','1','0','0','0','0','1','1','0','0'),
            ('1','1','1','0','1','1','0','0','0','0','1','1','1','0'),
            ('1','1','1','0','1','1','0','0','0','1','0','0','0','0'),
            ('1','1','1','0','1','1','0','0','0','1','0','0','1','0'),
            ('1','1','1','0','1','1','0','0','0','1','0','1','0','0'),
            ('1','1','1','0','1','1','0','0','0','1','0','1','1','0'),
            ('1','1','1','0','1','1','0','0','0','1','1','0','0','0'),
            ('1','1','1','0','1','1','0','0','0','1','1','0','1','0'),
            ('1','1','1','0','1','1','0','0','0','1','1','1','0','0'),
            ('1','1','1','0','1','1','0','0','0','1','1','1','1','0'),
            ('1','1','1','0','1','1','0','0','1','0','0','0','0','0'),
            ('1','1','1','0','1','1','0','0','1','0','0','0','1','0'),
            ('1','1','1','0','1','1','0','0','1','0','0','1','0','0'),
            ('1','1','1','0','1','1','0','0','1','0','0','1','1','0'),
            ('1','1','1','0','1','1','0','0','1','0','1','0','0','0'),
            ('1','1','1','0','1','1','0','0','1','0','1','0','1','0'),
            ('1','1','1','0','1','1','0','0','1','0','1','1','0','0'),
            ('1','1','1','0','1','1','0','0','1','0','1','1','1','0'),
            ('1','1','1','0','1','1','0','0','1','1','0','0','0','0'),
            ('1','1','1','0','1','1','0','0','1','1','0','0','1','0'),
            ('1','1','1','0','1','1','0','0','1','1','0','1','0','0'),
            ('1','1','1','0','1','1','0','0','1','1','0','1','1','0'),
            ('1','1','1','0','1','1','0','0','1','1','1','0','0','0'),
            ('1','1','1','0','1','1','0','0','1','1','1','0','1','0'),
            ('1','1','1','0','1','1','0','0','1','1','1','1','0','0'),
            ('1','1','1','0','1','1','0','0','1','1','1','1','1','0'),
            ('1','1','1','0','1','1','0','1','0','0','0','0','0','0'),
            ('1','1','1','0','1','1','0','1','0','0','0','0','1','0'),
            ('1','1','1','0','1','1','0','1','0','0','0','1','0','0'),
            ('1','1','1','0','1','1','0','1','0','0','0','1','1','0'),
            ('1','1','1','0','1','1','0','1','0','0','1','0','0','0'),
            ('1','1','1','0','1','1','0','1','0','0','1','0','1','0'),
            ('1','1','1','0','1','1','0','1','0','0','1','1','0','0'),
            ('1','1','1','0','1','1','0','1','0','0','1','1','1','0'),
            ('1','1','1','0','1','1','0','1','0','1','0','0','0','0'),
            ('1','1','1','0','1','1','0','1','0','1','0','0','1','0'),
            ('1','1','1','0','1','1','0','1','0','1','0','1','0','0'),
            ('1','1','1','0','1','1','0','1','0','1','0','1','1','0'),
            ('1','1','1','0','1','1','0','1','0','1','1','0','0','0'),
            ('1','1','1','0','1','1','0','1','0','1','1','0','1','0'),
            ('1','1','1','0','1','1','0','1','0','1','1','1','0','0'),
            ('1','1','1','0','1','1','0','1','0','1','1','1','1','0'),
            ('1','1','1','0','1','1','0','1','1','0','0','0','0','0'),
            ('1','1','1','0','1','1','0','1','1','0','0','0','1','0'),
            ('1','1','1','0','1','1','0','1','1','0','0','1','0','0'),
            ('1','1','1','0','1','1','0','1','1','0','0','1','1','0'),
            ('1','1','1','0','1','1','0','1','1','0','1','0','0','0'),
            ('1','1','1','0','1','1','0','1','1','0','1','0','1','0'),
            ('1','1','1','0','1','1','0','1','1','0','1','1','0','0'),
            ('1','1','1','0','1','1','0','1','1','0','1','1','1','0'),
            ('1','1','1','0','1','1','0','1','1','1','0','0','0','0'),
            ('1','1','1','0','1','1','0','1','1','1','0','0','1','0'),
            ('1','1','1','0','1','1','0','1','1','1','0','1','0','0'),
            ('1','1','1','0','1','1','0','1','1','1','0','1','1','0'),
            ('1','1','1','0','1','1','0','1','1','1','1','0','0','0'),
            ('1','1','1','0','1','1','0','1','1','1','1','0','1','0'),
            ('1','1','1','0','1','1','0','1','1','1','1','1','0','0'),
            ('1','1','1','0','1','1','0','1','1','1','1','1','1','0'),
            ('1','1','1','0','1','1','1','0','0','0','0','0','0','0'),
            ('1','1','1','0','1','1','1','0','0','0','0','0','1','0'),
            ('1','1','1','0','1','1','1','0','0','0','0','1','0','0'),
            ('1','1','1','0','1','1','1','0','0','0','0','1','1','0'),
            ('1','1','1','0','1','1','1','0','0','0','1','0','0','0'),
            ('1','1','1','0','1','1','1','0','0','0','1','0','1','0'),
            ('1','1','1','0','1','1','1','0','0','0','1','1','0','0'),
            ('1','1','1','0','1','1','1','0','0','0','1','1','1','0'),
            ('1','1','1','0','1','1','1','0','0','1','0','0','0','0'),
            ('1','1','1','0','1','1','1','0','0','1','0','0','1','0'),
            ('1','1','1','0','1','1','1','0','0','1','0','1','0','0'),
            ('1','1','1','0','1','1','1','0','0','1','0','1','1','0'),
            ('1','1','1','0','1','1','1','0','0','1','1','0','0','0'),
            ('1','1','1','0','1','1','1','0','0','1','1','0','1','0'),
            ('1','1','1','0','1','1','1','0','0','1','1','1','0','0'),
            ('1','1','1','0','1','1','1','0','0','1','1','1','1','0'),
            ('1','1','1','0','1','1','1','0','1','0','0','0','0','0'),
            ('1','1','1','0','1','1','1','0','1','0','0','0','1','0'),
            ('1','1','1','0','1','1','1','0','1','0','0','1','0','0'),
            ('1','1','1','0','1','1','1','0','1','0','0','1','1','0'),
            ('1','1','1','0','1','1','1','0','1','0','1','0','0','0'),
            ('1','1','1','0','1','1','1','0','1','0','1','0','1','0'),
            ('1','1','1','0','1','1','1','0','1','0','1','1','0','0'),
            ('1','1','1','0','1','1','1','0','1','0','1','1','1','0'),
            ('1','1','1','0','1','1','1','0','1','1','0','0','0','0'),
            ('1','1','1','0','1','1','1','0','1','1','0','0','1','0'),
            ('1','1','1','0','1','1','1','0','1','1','0','1','0','0'),
            ('1','1','1','0','1','1','1','0','1','1','0','1','1','0'),
            ('1','1','1','0','1','1','1','0','1','1','1','0','0','0'),
            ('1','1','1','0','1','1','1','0','1','1','1','0','1','0'),
            ('1','1','1','0','1','1','1','0','1','1','1','1','0','0'),
            ('1','1','1','0','1','1','1','0','1','1','1','1','1','0'),
            ('1','1','1','0','1','1','1','1','0','0','0','0','0','0'),
            ('1','1','1','0','1','1','1','1','0','0','0','0','1','0'),
            ('1','1','1','0','1','1','1','1','0','0','0','1','0','0'),
            ('1','1','1','0','1','1','1','1','0','0','0','1','1','0'),
            ('1','1','1','0','1','1','1','1','0','0','1','0','0','0'),
            ('1','1','1','0','1','1','1','1','0','0','1','0','1','0'),
            ('1','1','1','0','1','1','1','1','0','0','1','1','0','0'),
            ('1','1','1','0','1','1','1','1','0','0','1','1','1','0'),
            ('1','1','1','0','1','1','1','1','0','1','0','0','0','0'),
            ('1','1','1','0','1','1','1','1','0','1','0','0','1','0'),
            ('1','1','1','0','1','1','1','1','0','1','0','1','0','0'),
            ('1','1','1','0','1','1','1','1','0','1','0','1','1','0'),
            ('1','1','1','0','1','1','1','1','0','1','1','0','0','0'),
            ('1','1','1','0','1','1','1','1','0','1','1','0','1','0'),
            ('1','1','1','0','1','1','1','1','0','1','1','1','0','0'),
            ('1','1','1','0','1','1','1','1','0','1','1','1','1','0'),
            ('1','1','1','0','1','1','1','1','1','0','0','0','0','0'),
            ('1','1','1','0','1','1','1','1','1','0','0','0','1','0'),
            ('1','1','1','0','1','1','1','1','1','0','0','1','0','0'),
            ('1','1','1','0','1','1','1','1','1','0','0','1','1','0'),
            ('1','1','1','0','1','1','1','1','1','0','1','0','0','0'),
            ('1','1','1','0','1','1','1','1','1','0','1','0','1','0'),
            ('1','1','1','0','1','1','1','1','1','0','1','1','0','0'),
            ('1','1','1','0','1','1','1','1','1','0','1','1','1','0'),
            ('1','1','1','0','1','1','1','1','1','1','0','0','0','0'),
            ('1','1','1','0','1','1','1','1','1','1','0','0','1','0'),
            ('1','1','1','0','1','1','1','1','1','1','0','1','0','0'),
            ('1','1','1','0','1','1','1','1','1','1','0','1','1','0'),
            ('1','1','1','0','1','1','1','1','1','1','1','0','0','0'),
            ('1','1','1','0','1','1','1','1','1','1','1','0','1','0'),
            ('1','1','1','0','1','1','1','1','1','1','1','1','0','0'),
            ('1','1','1','0','1','1','1','1','1','1','1','1','1','0'),
            ('1','1','1','1','0','0','0','0','0','0','0','0','0','0'),
            ('1','1','1','1','0','0','0','0','0','0','0','0','1','0'),
            ('1','1','1','1','0','0','0','0','0','0','0','1','0','0'),
            ('1','1','1','1','0','0','0','0','0','0','0','1','1','0'),
            ('1','1','1','1','0','0','0','0','0','0','1','0','0','0'),
            ('1','1','1','1','0','0','0','0','0','0','1','0','1','0'),
            ('1','1','1','1','0','0','0','0','0','0','1','1','0','0'),
            ('1','1','1','1','0','0','0','0','0','0','1','1','1','0'),
            ('1','1','1','1','0','0','0','0','0','1','0','0','0','0'),
            ('1','1','1','1','0','0','0','0','0','1','0','0','1','0'),
            ('1','1','1','1','0','0','0','0','0','1','0','1','0','0'),
            ('1','1','1','1','0','0','0','0','0','1','0','1','1','0'),
            ('1','1','1','1','0','0','0','0','0','1','1','0','0','0'),
            ('1','1','1','1','0','0','0','0','0','1','1','0','1','0'),
            ('1','1','1','1','0','0','0','0','0','1','1','1','0','0'),
            ('1','1','1','1','0','0','0','0','0','1','1','1','1','0'),
            ('1','1','1','1','0','0','0','0','1','0','0','0','0','0'),
            ('1','1','1','1','0','0','0','0','1','0','0','0','1','0'),
            ('1','1','1','1','0','0','0','0','1','0','0','1','0','0'),
            ('1','1','1','1','0','0','0','0','1','0','0','1','1','0'),
            ('1','1','1','1','0','0','0','0','1','0','1','0','0','0'),
            ('1','1','1','1','0','0','0','0','1','0','1','0','1','0'),
            ('1','1','1','1','0','0','0','0','1','0','1','1','0','0'),
            ('1','1','1','1','0','0','0','0','1','0','1','1','1','0'),
            ('1','1','1','1','0','0','0','0','1','1','0','0','0','0'),
            ('1','1','1','1','0','0','0','0','1','1','0','0','1','0'),
            ('1','1','1','1','0','0','0','0','1','1','0','1','0','0'),
            ('1','1','1','1','0','0','0','0','1','1','0','1','1','0'),
            ('1','1','1','1','0','0','0','0','1','1','1','0','0','0'),
            ('1','1','1','1','0','0','0','0','1','1','1','0','1','0'),
            ('1','1','1','1','0','0','0','0','1','1','1','1','0','0'),
            ('1','1','1','1','0','0','0','0','1','1','1','1','1','0'),
            ('1','1','1','1','0','0','0','1','0','0','0','0','0','0'),
            ('1','1','1','1','0','0','0','1','0','0','0','0','1','0'),
            ('1','1','1','1','0','0','0','1','0','0','0','1','0','0'),
            ('1','1','1','1','0','0','0','1','0','0','0','1','1','0'),
            ('1','1','1','1','0','0','0','1','0','0','1','0','0','0'),
            ('1','1','1','1','0','0','0','1','0','0','1','0','1','0'),
            ('1','1','1','1','0','0','0','1','0','0','1','1','0','0'),
            ('1','1','1','1','0','0','0','1','0','0','1','1','1','0'),
            ('1','1','1','1','0','0','0','1','0','1','0','0','0','0'),
            ('1','1','1','1','0','0','0','1','0','1','0','0','1','0'),
            ('1','1','1','1','0','0','0','1','0','1','0','1','0','0'),
            ('1','1','1','1','0','0','0','1','0','1','0','1','1','0'),
            ('1','1','1','1','0','0','0','1','0','1','1','0','0','0'),
            ('1','1','1','1','0','0','0','1','0','1','1','0','1','0'),
            ('1','1','1','1','0','0','0','1','0','1','1','1','0','0'),
            ('1','1','1','1','0','0','0','1','0','1','1','1','1','0'),
            ('1','1','1','1','0','0','0','1','1','0','0','0','0','0'),
            ('1','1','1','1','0','0','0','1','1','0','0','0','1','0'),
            ('1','1','1','1','0','0','0','1','1','0','0','1','0','0'),
            ('1','1','1','1','0','0','0','1','1','0','0','1','1','0'),
            ('1','1','1','1','0','0','0','1','1','0','1','0','0','0'),
            ('1','1','1','1','0','0','0','1','1','0','1','0','1','0'),
            ('1','1','1','1','0','0','0','1','1','0','1','1','0','0'),
            ('1','1','1','1','0','0','0','1','1','0','1','1','1','0'),
            ('1','1','1','1','0','0','0','1','1','1','0','0','0','0'),
            ('1','1','1','1','0','0','0','1','1','1','0','0','1','0'),
            ('1','1','1','1','0','0','0','1','1','1','0','1','0','0'),
            ('1','1','1','1','0','0','0','1','1','1','0','1','1','0'),
            ('1','1','1','1','0','0','0','1','1','1','1','0','0','0'),
            ('1','1','1','1','0','0','0','1','1','1','1','0','1','0'),
            ('1','1','1','1','0','0','0','1','1','1','1','1','0','0'),
            ('1','1','1','1','0','0','0','1','1','1','1','1','1','0'),
            ('1','1','1','1','0','0','1','0','0','0','0','0','0','0'),
            ('1','1','1','1','0','0','1','0','0','0','0','0','1','0'),
            ('1','1','1','1','0','0','1','0','0','0','0','1','0','0'),
            ('1','1','1','1','0','0','1','0','0','0','0','1','1','0'),
            ('1','1','1','1','0','0','1','0','0','0','1','0','0','0'),
            ('1','1','1','1','0','0','1','0','0','0','1','0','1','0'),
            ('1','1','1','1','0','0','1','0','0','0','1','1','0','0'),
            ('1','1','1','1','0','0','1','0','0','0','1','1','1','0'),
            ('1','1','1','1','0','0','1','0','0','1','0','0','0','0'),
            ('1','1','1','1','0','0','1','0','0','1','0','0','1','0'),
            ('1','1','1','1','0','0','1','0','0','1','0','1','0','0'),
            ('1','1','1','1','0','0','1','0','0','1','0','1','1','0'),
            ('1','1','1','1','0','0','1','0','0','1','1','0','0','0'),
            ('1','1','1','1','0','0','1','0','0','1','1','0','1','0'),
            ('1','1','1','1','0','0','1','0','0','1','1','1','0','0'),
            ('1','1','1','1','0','0','1','0','0','1','1','1','1','0'),
            ('1','1','1','1','0','0','1','0','1','0','0','0','0','0'),
            ('1','1','1','1','0','0','1','0','1','0','0','0','1','0'),
            ('1','1','1','1','0','0','1','0','1','0','0','1','0','0'),
            ('1','1','1','1','0','0','1','0','1','0','0','1','1','0'),
            ('1','1','1','1','0','0','1','0','1','0','1','0','0','0'),
            ('1','1','1','1','0','0','1','0','1','0','1','0','1','0'),
            ('1','1','1','1','0','0','1','0','1','0','1','1','0','0'),
            ('1','1','1','1','0','0','1','0','1','0','1','1','1','0'),
            ('1','1','1','1','0','0','1','0','1','1','0','0','0','0'),
            ('1','1','1','1','0','0','1','0','1','1','0','0','1','0'),
            ('1','1','1','1','0','0','1','0','1','1','0','1','0','0'),
            ('1','1','1','1','0','0','1','0','1','1','0','1','1','0'),
            ('1','1','1','1','0','0','1','0','1','1','1','0','0','0'),
            ('1','1','1','1','0','0','1','0','1','1','1','0','1','0'),
            ('1','1','1','1','0','0','1','0','1','1','1','1','0','0'),
            ('1','1','1','1','0','0','1','0','1','1','1','1','1','0'),
            ('1','1','1','1','0','0','1','1','0','0','0','0','0','0'),
            ('1','1','1','1','0','0','1','1','0','0','0','0','1','0'),
            ('1','1','1','1','0','0','1','1','0','0','0','1','0','0'),
            ('1','1','1','1','0','0','1','1','0','0','0','1','1','0'),
            ('1','1','1','1','0','0','1','1','0','0','1','0','0','0'),
            ('1','1','1','1','0','0','1','1','0','0','1','0','1','0'),
            ('1','1','1','1','0','0','1','1','0','0','1','1','0','0'),
            ('1','1','1','1','0','0','1','1','0','0','1','1','1','0'),
            ('1','1','1','1','0','0','1','1','0','1','0','0','0','0'),
            ('1','1','1','1','0','0','1','1','0','1','0','0','1','0'),
            ('1','1','1','1','0','0','1','1','0','1','0','1','0','0'),
            ('1','1','1','1','0','0','1','1','0','1','0','1','1','0'),
            ('1','1','1','1','0','0','1','1','0','1','1','0','0','0'),
            ('1','1','1','1','0','0','1','1','0','1','1','0','1','0'),
            ('1','1','1','1','0','0','1','1','0','1','1','1','0','0'),
            ('1','1','1','1','0','0','1','1','0','1','1','1','1','0'),
            ('1','1','1','1','0','0','1','1','1','0','0','0','0','0'),
            ('1','1','1','1','0','0','1','1','1','0','0','0','1','0'),
            ('1','1','1','1','0','0','1','1','1','0','0','1','0','0'),
            ('1','1','1','1','0','0','1','1','1','0','0','1','1','0'),
            ('1','1','1','1','0','0','1','1','1','0','1','0','0','0'),
            ('1','1','1','1','0','0','1','1','1','0','1','0','1','0'),
            ('1','1','1','1','0','0','1','1','1','0','1','1','0','0'),
            ('1','1','1','1','0','0','1','1','1','0','1','1','1','0'),
            ('1','1','1','1','0','0','1','1','1','1','0','0','0','0'),
            ('1','1','1','1','0','0','1','1','1','1','0','0','1','0'),
            ('1','1','1','1','0','0','1','1','1','1','0','1','0','0'),
            ('1','1','1','1','0','0','1','1','1','1','0','1','1','0'),
            ('1','1','1','1','0','0','1','1','1','1','1','0','0','0'),
            ('1','1','1','1','0','0','1','1','1','1','1','0','1','0'),
            ('1','1','1','1','0','0','1','1','1','1','1','1','0','0'),
            ('1','1','1','1','0','0','1','1','1','1','1','1','1','0'),
            ('1','1','1','1','0','1','0','0','0','0','0','0','0','0'),
            ('1','1','1','1','0','1','0','0','0','0','0','0','1','0'),
            ('1','1','1','1','0','1','0','0','0','0','0','1','0','0'),
            ('1','1','1','1','0','1','0','0','0','0','0','1','1','0'),
            ('1','1','1','1','0','1','0','0','0','0','1','0','0','0'),
            ('1','1','1','1','0','1','0','0','0','0','1','0','1','0'),
            ('1','1','1','1','0','1','0','0','0','0','1','1','0','0'),
            ('1','1','1','1','0','1','0','0','0','0','1','1','1','0'),
            ('1','1','1','1','0','1','0','0','0','1','0','0','0','0'),
            ('1','1','1','1','0','1','0','0','0','1','0','0','1','0'),
            ('1','1','1','1','0','1','0','0','0','1','0','1','0','0'),
            ('1','1','1','1','0','1','0','0','0','1','0','1','1','0'),
            ('1','1','1','1','0','1','0','0','0','1','1','0','0','0'),
            ('1','1','1','1','0','1','0','0','0','1','1','0','1','0'),
            ('1','1','1','1','0','1','0','0','0','1','1','1','0','0'),
            ('1','1','1','1','0','1','0','0','0','1','1','1','1','0'),
            ('1','1','1','1','0','1','0','0','1','0','0','0','0','0'),
            ('1','1','1','1','0','1','0','0','1','0','0','0','1','0'),
            ('1','1','1','1','0','1','0','0','1','0','0','1','0','0'),
            ('1','1','1','1','0','1','0','0','1','0','0','1','1','0'),
            ('1','1','1','1','0','1','0','0','1','0','1','0','0','0'),
            ('1','1','1','1','0','1','0','0','1','0','1','0','1','0'),
            ('1','1','1','1','0','1','0','0','1','0','1','1','0','0'),
            ('1','1','1','1','0','1','0','0','1','0','1','1','1','0'),
            ('1','1','1','1','0','1','0','0','1','1','0','0','0','0'),
            ('1','1','1','1','0','1','0','0','1','1','0','0','1','0'),
            ('1','1','1','1','0','1','0','0','1','1','0','1','0','0'),
            ('1','1','1','1','0','1','0','0','1','1','0','1','1','0'),
            ('1','1','1','1','0','1','0','0','1','1','1','0','0','0'),
            ('1','1','1','1','0','1','0','0','1','1','1','0','1','0'),
            ('1','1','1','1','0','1','0','0','1','1','1','1','0','0'),
            ('1','1','1','1','0','1','0','0','1','1','1','1','1','0'),
            ('1','1','1','1','0','1','0','1','0','0','0','0','0','0'),
            ('1','1','1','1','0','1','0','1','0','0','0','0','1','0'),
            ('1','1','1','1','0','1','0','1','0','0','0','1','0','0'),
            ('1','1','1','1','0','1','0','1','0','0','0','1','1','0'),
            ('1','1','1','1','0','1','0','1','0','0','1','0','0','0'),
            ('1','1','1','1','0','1','0','1','0','0','1','0','1','0'),
            ('1','1','1','1','0','1','0','1','0','0','1','1','0','0'),
            ('1','1','1','1','0','1','0','1','0','0','1','1','1','0'),
            ('1','1','1','1','0','1','0','1','0','1','0','0','0','0'),
            ('1','1','1','1','0','1','0','1','0','1','0','0','1','0'),
            ('1','1','1','1','0','1','0','1','0','1','0','1','0','0'),
            ('1','1','1','1','0','1','0','1','0','1','0','1','1','0'),
            ('1','1','1','1','0','1','0','1','0','1','1','0','0','0'),
            ('1','1','1','1','0','1','0','1','0','1','1','0','1','0'),
            ('1','1','1','1','0','1','0','1','0','1','1','1','0','0'),
            ('1','1','1','1','0','1','0','1','0','1','1','1','1','0'),
            ('1','1','1','1','0','1','0','1','1','0','0','0','0','0'),
            ('1','1','1','1','0','1','0','1','1','0','0','0','1','0'),
            ('1','1','1','1','0','1','0','1','1','0','0','1','0','0'),
            ('1','1','1','1','0','1','0','1','1','0','0','1','1','0'),
            ('1','1','1','1','0','1','0','1','1','0','1','0','0','0'),
            ('1','1','1','1','0','1','0','1','1','0','1','0','1','0'),
            ('1','1','1','1','0','1','0','1','1','0','1','1','0','0'),
            ('1','1','1','1','0','1','0','1','1','0','1','1','1','0'),
            ('1','1','1','1','0','1','0','1','1','1','0','0','0','0'),
            ('1','1','1','1','0','1','0','1','1','1','0','0','1','0'),
            ('1','1','1','1','0','1','0','1','1','1','0','1','0','0'),
            ('1','1','1','1','0','1','0','1','1','1','0','1','1','0'),
            ('1','1','1','1','0','1','0','1','1','1','1','0','0','0'),
            ('1','1','1','1','0','1','0','1','1','1','1','0','1','0'),
            ('1','1','1','1','0','1','0','1','1','1','1','1','0','0'),
            ('1','1','1','1','0','1','0','1','1','1','1','1','1','0'),
            ('1','1','1','1','0','1','1','0','0','0','0','0','0','0'),
            ('1','1','1','1','0','1','1','0','0','0','0','0','1','0'),
            ('1','1','1','1','0','1','1','0','0','0','0','1','0','0'),
            ('1','1','1','1','0','1','1','0','0','0','0','1','1','0'),
            ('1','1','1','1','0','1','1','0','0','0','1','0','0','0'),
            ('1','1','1','1','0','1','1','0','0','0','1','0','1','0'),
            ('1','1','1','1','0','1','1','0','0','0','1','1','0','0'),
            ('1','1','1','1','0','1','1','0','0','0','1','1','1','0'),
            ('1','1','1','1','0','1','1','0','0','1','0','0','0','0'),
            ('1','1','1','1','0','1','1','0','0','1','0','0','1','0'),
            ('1','1','1','1','0','1','1','0','0','1','0','1','0','0'),
            ('1','1','1','1','0','1','1','0','0','1','0','1','1','0'),
            ('1','1','1','1','0','1','1','0','0','1','1','0','0','0'),
            ('1','1','1','1','0','1','1','0','0','1','1','0','1','0'),
            ('1','1','1','1','0','1','1','0','0','1','1','1','0','0'),
            ('1','1','1','1','0','1','1','0','0','1','1','1','1','0'),
            ('1','1','1','1','0','1','1','0','1','0','0','0','0','0'),
            ('1','1','1','1','0','1','1','0','1','0','0','0','1','0'),
            ('1','1','1','1','0','1','1','0','1','0','0','1','0','0'),
            ('1','1','1','1','0','1','1','0','1','0','0','1','1','0'),
            ('1','1','1','1','0','1','1','0','1','0','1','0','0','0'),
            ('1','1','1','1','0','1','1','0','1','0','1','0','1','0'),
            ('1','1','1','1','0','1','1','0','1','0','1','1','0','0'),
            ('1','1','1','1','0','1','1','0','1','0','1','1','1','0'),
            ('1','1','1','1','0','1','1','0','1','1','0','0','0','0'),
            ('1','1','1','1','0','1','1','0','1','1','0','0','1','0'),
            ('1','1','1','1','0','1','1','0','1','1','0','1','0','0'),
            ('1','1','1','1','0','1','1','0','1','1','0','1','1','0'),
            ('1','1','1','1','0','1','1','0','1','1','1','0','0','0'),
            ('1','1','1','1','0','1','1','0','1','1','1','0','1','0'),
            ('1','1','1','1','0','1','1','0','1','1','1','1','0','0'),
            ('1','1','1','1','0','1','1','0','1','1','1','1','1','0'),
            ('1','1','1','1','0','1','1','1','0','0','0','0','0','0'),
            ('1','1','1','1','0','1','1','1','0','0','0','0','1','0'),
            ('1','1','1','1','0','1','1','1','0','0','0','1','0','0'),
            ('1','1','1','1','0','1','1','1','0','0','0','1','1','0'),
            ('1','1','1','1','0','1','1','1','0','0','1','0','0','0'),
            ('1','1','1','1','0','1','1','1','0','0','1','0','1','0'),
            ('1','1','1','1','0','1','1','1','0','0','1','1','0','0'),
            ('1','1','1','1','0','1','1','1','0','0','1','1','1','0'),
            ('1','1','1','1','0','1','1','1','0','1','0','0','0','0'),
            ('1','1','1','1','0','1','1','1','0','1','0','0','1','0'),
            ('1','1','1','1','0','1','1','1','0','1','0','1','0','0'),
            ('1','1','1','1','0','1','1','1','0','1','0','1','1','0'),
            ('1','1','1','1','0','1','1','1','0','1','1','0','0','0'),
            ('1','1','1','1','0','1','1','1','0','1','1','0','1','0'),
            ('1','1','1','1','0','1','1','1','0','1','1','1','0','0'),
            ('1','1','1','1','0','1','1','1','0','1','1','1','1','0'),
            ('1','1','1','1','0','1','1','1','1','0','0','0','0','0'),
            ('1','1','1','1','0','1','1','1','1','0','0','0','1','0'),
            ('1','1','1','1','0','1','1','1','1','0','0','1','0','0'),
            ('1','1','1','1','0','1','1','1','1','0','0','1','1','0'),
            ('1','1','1','1','0','1','1','1','1','0','1','0','0','0'),
            ('1','1','1','1','0','1','1','1','1','0','1','0','1','0'),
            ('1','1','1','1','0','1','1','1','1','0','1','1','0','0'),
            ('1','1','1','1','0','1','1','1','1','0','1','1','1','0'),
            ('1','1','1','1','0','1','1','1','1','1','0','0','0','0'),
            ('1','1','1','1','0','1','1','1','1','1','0','0','1','0'),
            ('1','1','1','1','0','1','1','1','1','1','0','1','0','0'),
            ('1','1','1','1','0','1','1','1','1','1','0','1','1','0'),
            ('1','1','1','1','0','1','1','1','1','1','1','0','0','0'),
            ('1','1','1','1','0','1','1','1','1','1','1','0','1','0'),
            ('1','1','1','1','0','1','1','1','1','1','1','1','0','0'),
            ('1','1','1','1','0','1','1','1','1','1','1','1','1','0'),
            ('1','1','1','1','1','0','0','0','0','0','0','0','0','0'),
            ('1','1','1','1','1','0','0','0','0','0','0','0','1','0'),
            ('1','1','1','1','1','0','0','0','0','0','0','1','0','0'),
            ('1','1','1','1','1','0','0','0','0','0','0','1','1','0'),
            ('1','1','1','1','1','0','0','0','0','0','1','0','0','0'),
            ('1','1','1','1','1','0','0','0','0','0','1','0','1','0'),
            ('1','1','1','1','1','0','0','0','0','0','1','1','0','0'),
            ('1','1','1','1','1','0','0','0','0','0','1','1','1','0'),
            ('1','1','1','1','1','0','0','0','0','1','0','0','0','0'),
            ('1','1','1','1','1','0','0','0','0','1','0','0','1','0'),
            ('1','1','1','1','1','0','0','0','0','1','0','1','0','0'),
            ('1','1','1','1','1','0','0','0','0','1','0','1','1','0'),
            ('1','1','1','1','1','0','0','0','0','1','1','0','0','0'),
            ('1','1','1','1','1','0','0','0','0','1','1','0','1','0'),
            ('1','1','1','1','1','0','0','0','0','1','1','1','0','0'),
            ('1','1','1','1','1','0','0','0','0','1','1','1','1','0'),
            ('1','1','1','1','1','0','0','0','1','0','0','0','0','0'),
            ('1','1','1','1','1','0','0','0','1','0','0','0','1','0'),
            ('1','1','1','1','1','0','0','0','1','0','0','1','0','0'),
            ('1','1','1','1','1','0','0','0','1','0','0','1','1','0'),
            ('1','1','1','1','1','0','0','0','1','0','1','0','0','0'),
            ('1','1','1','1','1','0','0','0','1','0','1','0','1','0'),
            ('1','1','1','1','1','0','0','0','1','0','1','1','0','0'),
            ('1','1','1','1','1','0','0','0','1','0','1','1','1','0'),
            ('1','1','1','1','1','0','0','0','1','1','0','0','0','0'),
            ('1','1','1','1','1','0','0','0','1','1','0','0','1','0'),
            ('1','1','1','1','1','0','0','0','1','1','0','1','0','0'),
            ('1','1','1','1','1','0','0','0','1','1','0','1','1','0'),
            ('1','1','1','1','1','0','0','0','1','1','1','0','0','0'),
            ('1','1','1','1','1','0','0','0','1','1','1','0','1','0'),
            ('1','1','1','1','1','0','0','0','1','1','1','1','0','0'),
            ('1','1','1','1','1','0','0','0','1','1','1','1','1','0'),
            ('1','1','1','1','1','0','0','1','0','0','0','0','0','0'),
            ('1','1','1','1','1','0','0','1','0','0','0','0','1','0'),
            ('1','1','1','1','1','0','0','1','0','0','0','1','0','0'),
            ('1','1','1','1','1','0','0','1','0','0','0','1','1','0'),
            ('1','1','1','1','1','0','0','1','0','0','1','0','0','0'),
            ('1','1','1','1','1','0','0','1','0','0','1','0','1','0'),
            ('1','1','1','1','1','0','0','1','0','0','1','1','0','0'),
            ('1','1','1','1','1','0','0','1','0','0','1','1','1','0'),
            ('1','1','1','1','1','0','0','1','0','1','0','0','0','0'),
            ('1','1','1','1','1','0','0','1','0','1','0','0','1','0'),
            ('1','1','1','1','1','0','0','1','0','1','0','1','0','0'),
            ('1','1','1','1','1','0','0','1','0','1','0','1','1','0'),
            ('1','1','1','1','1','0','0','1','0','1','1','0','0','0'),
            ('1','1','1','1','1','0','0','1','0','1','1','0','1','0'),
            ('1','1','1','1','1','0','0','1','0','1','1','1','0','0'),
            ('1','1','1','1','1','0','0','1','0','1','1','1','1','0'),
            ('1','1','1','1','1','0','0','1','1','0','0','0','0','0'),
            ('1','1','1','1','1','0','0','1','1','0','0','0','1','0'),
            ('1','1','1','1','1','0','0','1','1','0','0','1','0','0'),
            ('1','1','1','1','1','0','0','1','1','0','0','1','1','0'),
            ('1','1','1','1','1','0','0','1','1','0','1','0','0','0'),
            ('1','1','1','1','1','0','0','1','1','0','1','0','1','0'),
            ('1','1','1','1','1','0','0','1','1','0','1','1','0','0'),
            ('1','1','1','1','1','0','0','1','1','0','1','1','1','0'),
            ('1','1','1','1','1','0','0','1','1','1','0','0','0','0'),
            ('1','1','1','1','1','0','0','1','1','1','0','0','1','0'),
            ('1','1','1','1','1','0','0','1','1','1','0','1','0','0'),
            ('1','1','1','1','1','0','0','1','1','1','0','1','1','0'),
            ('1','1','1','1','1','0','0','1','1','1','1','0','0','0'),
            ('1','1','1','1','1','0','0','1','1','1','1','0','1','0'),
            ('1','1','1','1','1','0','0','1','1','1','1','1','0','0'),
            ('1','1','1','1','1','0','0','1','1','1','1','1','1','0'),
            ('1','1','1','1','1','0','1','0','0','0','0','0','0','0'),
            ('1','1','1','1','1','0','1','0','0','0','0','0','1','0'),
            ('1','1','1','1','1','0','1','0','0','0','0','1','0','0'),
            ('1','1','1','1','1','0','1','0','0','0','0','1','1','0'),
            ('1','1','1','1','1','0','1','0','0','0','1','0','0','0'),
            ('1','1','1','1','1','0','1','0','0','0','1','0','1','0'),
            ('1','1','1','1','1','0','1','0','0','0','1','1','0','0'),
            ('1','1','1','1','1','0','1','0','0','0','1','1','1','0'),
            ('1','1','1','1','1','0','1','0','0','1','0','0','0','0'),
            ('1','1','1','1','1','0','1','0','0','1','0','0','1','0'),
            ('1','1','1','1','1','0','1','0','0','1','0','1','0','0'),
            ('1','1','1','1','1','0','1','0','0','1','0','1','1','0'),
            ('1','1','1','1','1','0','1','0','0','1','1','0','0','0'),
            ('1','1','1','1','1','0','1','0','0','1','1','0','1','0'),
            ('1','1','1','1','1','0','1','0','0','1','1','1','0','0'),
            ('1','1','1','1','1','0','1','0','0','1','1','1','1','0'),
            ('1','1','1','1','1','0','1','0','1','0','0','0','0','0'),
            ('1','1','1','1','1','0','1','0','1','0','0','0','1','0'),
            ('1','1','1','1','1','0','1','0','1','0','0','1','0','0'),
            ('1','1','1','1','1','0','1','0','1','0','0','1','1','0'),
            ('1','1','1','1','1','0','1','0','1','0','1','0','0','0'),
            ('1','1','1','1','1','0','1','0','1','0','1','0','1','0'),
            ('1','1','1','1','1','0','1','0','1','0','1','1','0','0'),
            ('1','1','1','1','1','0','1','0','1','0','1','1','1','0'),
            ('1','1','1','1','1','0','1','0','1','1','0','0','0','0'),
            ('1','1','1','1','1','0','1','0','1','1','0','0','1','0'),
            ('1','1','1','1','1','0','1','0','1','1','0','1','0','0'),
            ('1','1','1','1','1','0','1','0','1','1','0','1','1','0'),
            ('1','1','1','1','1','0','1','0','1','1','1','0','0','0'),
            ('1','1','1','1','1','0','1','0','1','1','1','0','1','0'),
            ('1','1','1','1','1','0','1','0','1','1','1','1','0','0'),
            ('1','1','1','1','1','0','1','0','1','1','1','1','1','0'),
            ('1','1','1','1','1','0','1','1','0','0','0','0','0','0'),
            ('1','1','1','1','1','0','1','1','0','0','0','0','1','0'),
            ('1','1','1','1','1','0','1','1','0','0','0','1','0','0'),
            ('1','1','1','1','1','0','1','1','0','0','0','1','1','0'),
            ('1','1','1','1','1','0','1','1','0','0','1','0','0','0'),
            ('1','1','1','1','1','0','1','1','0','0','1','0','1','0'),
            ('1','1','1','1','1','0','1','1','0','0','1','1','0','0'),
            ('1','1','1','1','1','0','1','1','0','0','1','1','1','0'),
            ('1','1','1','1','1','0','1','1','0','1','0','0','0','0'),
            ('1','1','1','1','1','0','1','1','0','1','0','0','1','0'),
            ('1','1','1','1','1','0','1','1','0','1','0','1','0','0'),
            ('1','1','1','1','1','0','1','1','0','1','0','1','1','0'),
            ('1','1','1','1','1','0','1','1','0','1','1','0','0','0'),
            ('1','1','1','1','1','0','1','1','0','1','1','0','1','0'),
            ('1','1','1','1','1','0','1','1','0','1','1','1','0','0'),
            ('1','1','1','1','1','0','1','1','0','1','1','1','1','0'),
            ('1','1','1','1','1','0','1','1','1','0','0','0','0','0'),
            ('1','1','1','1','1','0','1','1','1','0','0','0','1','0'),
            ('1','1','1','1','1','0','1','1','1','0','0','1','0','0'),
            ('1','1','1','1','1','0','1','1','1','0','0','1','1','0'),
            ('1','1','1','1','1','0','1','1','1','0','1','0','0','0'),
            ('1','1','1','1','1','0','1','1','1','0','1','0','1','0'),
            ('1','1','1','1','1','0','1','1','1','0','1','1','0','0'),
            ('1','1','1','1','1','0','1','1','1','0','1','1','1','0'),
            ('1','1','1','1','1','0','1','1','1','1','0','0','0','0'),
            ('1','1','1','1','1','0','1','1','1','1','0','0','1','0'),
            ('1','1','1','1','1','0','1','1','1','1','0','1','0','0'),
            ('1','1','1','1','1','0','1','1','1','1','0','1','1','0'),
            ('1','1','1','1','1','0','1','1','1','1','1','0','0','0'),
            ('1','1','1','1','1','0','1','1','1','1','1','0','1','0'),
            ('1','1','1','1','1','0','1','1','1','1','1','1','0','0'),
            ('1','1','1','1','1','0','1','1','1','1','1','1','1','0'),
            ('1','1','1','1','1','1','0','0','0','0','0','0','0','0'),
            ('1','1','1','1','1','1','0','0','0','0','0','0','1','0'),
            ('1','1','1','1','1','1','0','0','0','0','0','1','0','0'),
            ('1','1','1','1','1','1','0','0','0','0','0','1','1','0'),
            ('1','1','1','1','1','1','0','0','0','0','1','0','0','0'),
            ('1','1','1','1','1','1','0','0','0','0','1','0','1','0'),
            ('1','1','1','1','1','1','0','0','0','0','1','1','0','0'),
            ('1','1','1','1','1','1','0','0','0','0','1','1','1','0'),
            ('1','1','1','1','1','1','0','0','0','1','0','0','0','0'),
            ('1','1','1','1','1','1','0','0','0','1','0','0','1','0'),
            ('1','1','1','1','1','1','0','0','0','1','0','1','0','0'),
            ('1','1','1','1','1','1','0','0','0','1','0','1','1','0'),
            ('1','1','1','1','1','1','0','0','0','1','1','0','0','0'),
            ('1','1','1','1','1','1','0','0','0','1','1','0','1','0'),
            ('1','1','1','1','1','1','0','0','0','1','1','1','0','0'),
            ('1','1','1','1','1','1','0','0','0','1','1','1','1','0'),
            ('1','1','1','1','1','1','0','0','1','0','0','0','0','0'),
            ('1','1','1','1','1','1','0','0','1','0','0','0','1','0'),
            ('1','1','1','1','1','1','0','0','1','0','0','1','0','0'),
            ('1','1','1','1','1','1','0','0','1','0','0','1','1','0'),
            ('1','1','1','1','1','1','0','0','1','0','1','0','0','0'),
            ('1','1','1','1','1','1','0','0','1','0','1','0','1','0'),
            ('1','1','1','1','1','1','0','0','1','0','1','1','0','0'),
            ('1','1','1','1','1','1','0','0','1','0','1','1','1','0'),
            ('1','1','1','1','1','1','0','0','1','1','0','0','0','0'),
            ('1','1','1','1','1','1','0','0','1','1','0','0','1','0'),
            ('1','1','1','1','1','1','0','0','1','1','0','1','0','0'),
            ('1','1','1','1','1','1','0','0','1','1','0','1','1','0'),
            ('1','1','1','1','1','1','0','0','1','1','1','0','0','0'),
            ('1','1','1','1','1','1','0','0','1','1','1','0','1','0'),
            ('1','1','1','1','1','1','0','0','1','1','1','1','0','0'),
            ('1','1','1','1','1','1','0','0','1','1','1','1','1','0'),
            ('1','1','1','1','1','1','0','1','0','0','0','0','0','0'),
            ('1','1','1','1','1','1','0','1','0','0','0','0','1','0'),
            ('1','1','1','1','1','1','0','1','0','0','0','1','0','0'),
            ('1','1','1','1','1','1','0','1','0','0','0','1','1','0'),
            ('1','1','1','1','1','1','0','1','0','0','1','0','0','0'),
            ('1','1','1','1','1','1','0','1','0','0','1','0','1','0'),
            ('1','1','1','1','1','1','0','1','0','0','1','1','0','0'),
            ('1','1','1','1','1','1','0','1','0','0','1','1','1','0'),
            ('1','1','1','1','1','1','0','1','0','1','0','0','0','0'),
            ('1','1','1','1','1','1','0','1','0','1','0','0','1','0'),
            ('1','1','1','1','1','1','0','1','0','1','0','1','0','0'),
            ('1','1','1','1','1','1','0','1','0','1','0','1','1','0'),
            ('1','1','1','1','1','1','0','1','0','1','1','0','0','0'),
            ('1','1','1','1','1','1','0','1','0','1','1','0','1','0'),
            ('1','1','1','1','1','1','0','1','0','1','1','1','0','0'),
            ('1','1','1','1','1','1','0','1','0','1','1','1','1','0'),
            ('1','1','1','1','1','1','0','1','1','0','0','0','0','0'),
            ('1','1','1','1','1','1','0','1','1','0','0','0','1','0'),
            ('1','1','1','1','1','1','0','1','1','0','0','1','0','0'),
            ('1','1','1','1','1','1','0','1','1','0','0','1','1','0'),
            ('1','1','1','1','1','1','0','1','1','0','1','0','0','0'),
            ('1','1','1','1','1','1','0','1','1','0','1','0','1','0'),
            ('1','1','1','1','1','1','0','1','1','0','1','1','0','0'),
            ('1','1','1','1','1','1','0','1','1','0','1','1','1','0'),
            ('1','1','1','1','1','1','0','1','1','1','0','0','0','0'),
            ('1','1','1','1','1','1','0','1','1','1','0','0','1','0'),
            ('1','1','1','1','1','1','0','1','1','1','0','1','0','0'),
            ('1','1','1','1','1','1','0','1','1','1','0','1','1','0'),
            ('1','1','1','1','1','1','0','1','1','1','1','0','0','0'),
            ('1','1','1','1','1','1','0','1','1','1','1','0','1','0'),
            ('1','1','1','1','1','1','0','1','1','1','1','1','0','0'),
            ('1','1','1','1','1','1','0','1','1','1','1','1','1','0'),
            ('1','1','1','1','1','1','1','0','0','0','0','0','0','0'),
            ('1','1','1','1','1','1','1','0','0','0','0','0','1','0'),
            ('1','1','1','1','1','1','1','0','0','0','0','1','0','0'),
            ('1','1','1','1','1','1','1','0','0','0','0','1','1','0'),
            ('1','1','1','1','1','1','1','0','0','0','1','0','0','0'),
            ('1','1','1','1','1','1','1','0','0','0','1','0','1','0'),
            ('1','1','1','1','1','1','1','0','0','0','1','1','0','0'),
            ('1','1','1','1','1','1','1','0','0','0','1','1','1','0'),
            ('1','1','1','1','1','1','1','0','0','1','0','0','0','0'),
            ('1','1','1','1','1','1','1','0','0','1','0','0','1','0'),
            ('1','1','1','1','1','1','1','0','0','1','0','1','0','0'),
            ('1','1','1','1','1','1','1','0','0','1','0','1','1','0'),
            ('1','1','1','1','1','1','1','0','0','1','1','0','0','0'),
            ('1','1','1','1','1','1','1','0','0','1','1','0','1','0'),
            ('1','1','1','1','1','1','1','0','0','1','1','1','0','0'),
            ('1','1','1','1','1','1','1','0','0','1','1','1','1','0'),
            ('1','1','1','1','1','1','1','0','1','0','0','0','0','0'),
            ('1','1','1','1','1','1','1','0','1','0','0','0','1','0'),
            ('1','1','1','1','1','1','1','0','1','0','0','1','0','0'),
            ('1','1','1','1','1','1','1','0','1','0','0','1','1','0'),
            ('1','1','1','1','1','1','1','0','1','0','1','0','0','0'),
            ('1','1','1','1','1','1','1','0','1','0','1','0','1','0'),
            ('1','1','1','1','1','1','1','0','1','0','1','1','0','0'),
            ('1','1','1','1','1','1','1','0','1','0','1','1','1','0'),
            ('1','1','1','1','1','1','1','0','1','1','0','0','0','0'),
            ('1','1','1','1','1','1','1','0','1','1','0','0','1','0'),
            ('1','1','1','1','1','1','1','0','1','1','0','1','0','0'),
            ('1','1','1','1','1','1','1','0','1','1','0','1','1','0'),
            ('1','1','1','1','1','1','1','0','1','1','1','0','0','0'),
            ('1','1','1','1','1','1','1','0','1','1','1','0','1','0'),
            ('1','1','1','1','1','1','1','0','1','1','1','1','0','0'),
            ('1','1','1','1','1','1','1','0','1','1','1','1','1','0'),
            ('1','1','1','1','1','1','1','1','0','0','0','0','0','0'),
            ('1','1','1','1','1','1','1','1','0','0','0','0','1','0'),
            ('1','1','1','1','1','1','1','1','0','0','0','1','0','0'),
            ('1','1','1','1','1','1','1','1','0','0','0','1','1','0'),
            ('1','1','1','1','1','1','1','1','0','0','1','0','0','0'),
            ('1','1','1','1','1','1','1','1','0','0','1','0','1','0'),
            ('1','1','1','1','1','1','1','1','0','0','1','1','0','0'),
            ('1','1','1','1','1','1','1','1','0','0','1','1','1','0'),
            ('1','1','1','1','1','1','1','1','0','1','0','0','0','0'),
            ('1','1','1','1','1','1','1','1','0','1','0','0','1','0'),
            ('1','1','1','1','1','1','1','1','0','1','0','1','0','0'),
            ('1','1','1','1','1','1','1','1','0','1','0','1','1','0'),
            ('1','1','1','1','1','1','1','1','0','1','1','0','0','0'),
            ('1','1','1','1','1','1','1','1','0','1','1','0','1','0'),
            ('1','1','1','1','1','1','1','1','0','1','1','1','0','0'),
            ('1','1','1','1','1','1','1','1','0','1','1','1','1','0'),
            ('1','1','1','1','1','1','1','1','1','0','0','0','0','0'),
            ('1','1','1','1','1','1','1','1','1','0','0','0','1','0'),
            ('1','1','1','1','1','1','1','1','1','0','0','1','0','0'),
            ('1','1','1','1','1','1','1','1','1','0','0','1','1','0'),
            ('1','1','1','1','1','1','1','1','1','0','1','0','0','0'),
            ('1','1','1','1','1','1','1','1','1','0','1','0','1','0'),
            ('1','1','1','1','1','1','1','1','1','0','1','1','0','0'),
            ('1','1','1','1','1','1','1','1','1','0','1','1','1','0'),
            ('1','1','1','1','1','1','1','1','1','1','0','0','0','0'),
            ('1','1','1','1','1','1','1','1','1','1','0','0','1','0'),
            ('1','1','1','1','1','1','1','1','1','1','0','1','0','0'),
            ('1','1','1','1','1','1','1','1','1','1','0','1','1','0'),
            ('1','1','1','1','1','1','1','1','1','1','1','0','0','0'),
            ('1','1','1','1','1','1','1','1','1','1','1','0','1','0'),
            ('1','1','1','1','1','1','1','1','1','1','1','1','0','0'),
            ('1','1','1','1','1','1','1','1','1','1','1','1','1','0')
            
            );
        begin
           for i in tabela_verdade'range loop
                d0 <= tabela_verdade(i).d0;
                d1 <= tabela_verdade(i).d1;
                d2 <= tabela_verdade(i).d2;
                d3 <= tabela_verdade(i).d3;
                d4 <= tabela_verdade(i).d4;
                d5 <= tabela_verdade(i).d5;
                d6 <= tabela_verdade(i).d6;
                d7 <= tabela_verdade(i).d7;
                c1 <= tabela_verdade(i).c1;
                c2 <= tabela_verdade(i).c2;
                c3 <= tabela_verdade(i).c3;
                c4 <= tabela_verdade(i).c4;
                c5 <= tabela_verdade(i).c5;
            wait for 1 ns;
        end loop;
            report "Fim teste";
            wait;
    end process estimulo_checagem;
end;