library ieee;
use ieee.std_logic_1164.all;

entity fulladder4 is
    port(
        A, B: in std_logic_vector(3 downto 0);
        CIN: in std_logic;
        S: out std_logic_vector(3 downto 0);
        COUT: out std_logic
    );
end entity;

architecture structural of fulladder4 is

-- SEU CODIGO AQUI

begin

-- SEU CODIGO AQUI
--
-- Voce DEVE escrever uma arquitetura estrutural.
-- Ou seja, DEVE instanciar as entidades fulladder1 e
-- interliga-las de forma a produzir um somador 
-- completo de 4 bits.

end architecture;
