library ieee;
use ieee.std_logic_1164.all;


entity teste is
    generic (
        N: natural := 3
    );
end entity;

architecture rtl of teste is
    signal sensors: std_logic_vector(0 to N-1);
    signal key, clock, siren : std_logic;
begin

    alarme_0: entity work.alarm(behavioral)
    generic map (N)
    port map (sensors => sensors,key => key, clock => clock, siren => siren);
    
    barulho: process is
        type strutura is record
            sensors: std_logic_vector(0 to N-1);
            key, clock, siren : std_logic;
        end record;
        type vet_alarme is array (natural range<>) of strutura;
        constant tabela : vet_alarme := 
        (
        --     s    k   c   si
            ("000",'0','0','0'),
            ("000",'1','1','0'),
            ("000",'1','0','0'),
            ("000",'1','1','0'),
            ("000",'1','0','0'),
            ("000",'1','1','0'),
            ("000",'1','0','0'),
            ("000",'1','1','0'),
            ("000",'1','0','0'),
            ("000",'1','1','0'),
            ("000",'1','0','0'),
            ("000",'1','1','0'),
            ("000",'1','0','0'),
            ("000",'1','1','0'),
            ("000",'1','0','0'),
            ("000",'1','1','0'),
            ("000",'1','0','0'),
            ("000",'1','1','0'),
            ("000",'1','0','0'),
            ("000",'1','1','0'),
            ("000",'1','0','0'),
            ("000",'1','1','0'),
            ("000",'1','0','0'),
            ("000",'1','1','0'),
            ("000",'1','0','0'),
            ("000",'1','1','0'),
            ("000",'1','0','0'),
            ("000",'1','1','0'),
            ("000",'1','0','0'),
            ("000",'1','1','0'),
            ("000",'1','0','0'),
            ("000",'1','1','0'),
            ("000",'1','0','0'), 
            ("001",'1','1','0'), 
            ("001",'1','0','0'),
            ("001",'1','1','0'),
            ("001",'1','0','0'),
            ("001",'1','1','0'),
            ("001",'1','0','0'),
            ("001",'1','1','0'),
            ("001",'1','0','0'),
            ("001",'1','1','0'),
            ("001",'1','0','0'),
            ("001",'1','1','0'),
            ("001",'1','0','0'),
            ("001",'1','1','0'),
            ("001",'1','0','0'),
            ("001",'1','1','0'),
            ("001",'1','0','0'),
            ("001",'1','1','0'),
            ("001",'1','0','0'),
            ("001",'1','1','0'),
            ("001",'1','0','0'),
            ("010",'1','1','0'),
            ("010",'1','0','0'),
            ("010",'1','1','0'),
            ("010",'1','0','0'),
            ("010",'1','1','0'),
            ("100",'1','0','0'),
            ("100",'1','1','0'),
            ("100",'1','0','0'),
            ("100",'1','1','0'),
            ("100",'1','0','0'),
            ("100",'1','1','0'),
            ("100",'1','0','1'),
            ("100",'1','1','1'),
            ("100",'1','0','1'),
            ("100",'1','1','1'),
            ("000",'1','0','0'),
            ("000",'1','1','0'),
            ("000",'1','0','0'),
            ("000",'1','1','0'),
            ("000",'1','0','0'),
            ("000",'1','1','0'),
            ("000",'1','0','0'),
            ("000",'1','1','0'),
            ("000",'1','0','0'),
            ("000",'1','1','0'),
            ("000",'1','0','0'),
            ("000",'1','1','0'),
            ("000",'1','0','0'),
            ("000",'1','1','0'),
            ("000",'1','0','0'),
            ("000",'1','1','0'),
            ("000",'1','0','0'),
            ("000",'1','1','0'),
            ("000",'1','0','0'),
            ("000",'1','1','0'),
            ("000",'1','0','0'),
            ("000",'1','1','0'),
            ("000",'1','0','0'),
            ("000",'1','1','0'),
            ("000",'1','0','0'),
            ("000",'1','1','0'),
            ("000",'1','0','0'),
            ("000",'1','1','0'),
            ("000",'1','0','0'),
            ("000",'1','1','0'),
            ("000",'1','0','0'),
            ("000",'1','1','0'),
            ("000",'1','0','0'), 
            ("001",'1','1','0'), 
            ("001",'1','0','0'),
            ("001",'1','1','0'),
            ("001",'1','0','0'),
            ("001",'1','1','0'),
            ("001",'1','0','0'),
            ("001",'1','1','0'),
            ("001",'1','0','0'),
            ("001",'1','1','0'),
            ("001",'1','0','0'),
            ("001",'1','1','0'),
            ("001",'1','0','0'),
            ("001",'1','1','0'),
            ("001",'1','0','0'),
            ("001",'1','1','0'),
            ("001",'1','0','0'),
            ("001",'1','1','0'),
            ("001",'1','0','0'),
            ("001",'1','1','0'),
            ("001",'1','0','0'),
            ("010",'1','1','0'),
            ("010",'1','0','0'),
            ("010",'1','1','0'),
            ("010",'1','0','0'),
            ("010",'1','1','0'),
            ("100",'1','0','0'),
            ("100",'1','1','0'),
            ("100",'1','0','0'),
            ("100",'1','1','0'),
            ("100",'1','0','0'),
            ("100",'1','1','0'),
            ("100",'1','0','1'),
            ("100",'1','1','1'),
            ("100",'1','0','1'),
            ("100",'1','1','1')
        );
    begin
        for i in tabela'range loop
            sensors <= tabela(i).sensors;
            key <= tabela(i).key;
            clock <= tabela(i).clock;

            wait for 1 ns;

            assert siren = tabela(i).siren
                report "Sirene = " & std_logic'image(siren) &  " " & "No tempo = " & natural'image(i) 
                & " Era para ser = " & std_logic'image(tabela(i).siren);
        end loop;
            report "Fim processo!!!";
        wait;
    end process;
end architecture;